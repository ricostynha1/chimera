// This program was cloned from: https://github.com/Nilesh002/Multiplication-and-Accumulation-Unit-MAC-
// License: MIT License

module adder24(a,b,s);
input [23:0]a,b;
output [23:0]s;

assign s=a+b;

endmodule
