// This program was cloned from: https://github.com/thinkoco/de10-nano-riscv
// License: Apache License 2.0

//Created atTue Feb 19 16:05:10 2019
// This file created by ROM_V_Generator, a perl tool by DeeZeng

module BootROM(
  input clock,
  input oe,
  input me,
  input [10:0] address,
  output [31:0] q
);
  reg [31:0] out;
  reg [31:0] rom [0:2047];

  always @(posedge clock) begin
    if (me) begin
	  case(address)
             0:out <= 32'hf1402573;
             1:out <= 32'h00000597;
             2:out <= 32'h01058593;
             3:out <= 32'h200002b7;
             4:out <= 32'h00028067;
             5:out <= 32'hedfe0dd0;
             6:out <= 32'he80d0000;
             7:out <= 32'h38000000;
             8:out <= 32'h800c0000;
             9:out <= 32'h28000000;
             10:out <= 32'h11000000;
             11:out <= 32'h10000000;
             12:out <= 32'h00000000;
             13:out <= 32'h68010000;
             14:out <= 32'h480c0000;
             15:out <= 32'h00000000;
             16:out <= 32'h00000000;
             17:out <= 32'h00000000;
             18:out <= 32'h00000000;
             19:out <= 32'h01000000;
             20:out <= 32'h00000000;
             21:out <= 32'h03000000;
             22:out <= 32'h04000000;
             23:out <= 32'h00000000;
             24:out <= 32'h01000000;
             25:out <= 32'h03000000;
             26:out <= 32'h04000000;
             27:out <= 32'h0f000000;
             28:out <= 32'h01000000;
             29:out <= 32'h03000000;
             30:out <= 32'h21000000;
             31:out <= 32'h1b000000;
             32:out <= 32'h65657266;
             33:out <= 32'h70696863;
             34:out <= 32'h6f722c73;
             35:out <= 32'h74656b63;
             36:out <= 32'h70696863;
             37:out <= 32'h6b6e752d;
             38:out <= 32'h6e776f6e;
             39:out <= 32'h7665642d;
             40:out <= 32'h00000000;
             41:out <= 32'h03000000;
             42:out <= 32'h1d000000;
             43:out <= 32'h26000000;
             44:out <= 32'h65657266;
             45:out <= 32'h70696863;
             46:out <= 32'h6f722c73;
             47:out <= 32'h74656b63;
             48:out <= 32'h70696863;
             49:out <= 32'h6b6e752d;
             50:out <= 32'h6e776f6e;
             51:out <= 32'h00000000;
             52:out <= 32'h01000000;
             53:out <= 32'h61696c61;
             54:out <= 32'h00736573;
             55:out <= 32'h03000000;
             56:out <= 32'h15000000;
             57:out <= 32'h2c000000;
             58:out <= 32'h636f732f;
             59:out <= 32'h7265732f;
             60:out <= 32'h406c6169;
             61:out <= 32'h31303031;
             62:out <= 32'h30303033;
             63:out <= 32'h00000000;
             64:out <= 32'h03000000;
             65:out <= 32'h15000000;
             66:out <= 32'h34000000;
             67:out <= 32'h636f732f;
             68:out <= 32'h7265732f;
             69:out <= 32'h406c6169;
             70:out <= 32'h32303031;
             71:out <= 32'h30303033;
             72:out <= 32'h00000000;
             73:out <= 32'h02000000;
             74:out <= 32'h01000000;
             75:out <= 32'h73757063;
             76:out <= 32'h00000000;
             77:out <= 32'h03000000;
             78:out <= 32'h04000000;
             79:out <= 32'h00000000;
             80:out <= 32'h01000000;
             81:out <= 32'h03000000;
             82:out <= 32'h04000000;
             83:out <= 32'h0f000000;
             84:out <= 32'h00000000;
             85:out <= 32'h01000000;
             86:out <= 32'h40757063;
             87:out <= 32'h00000030;
             88:out <= 32'h03000000;
             89:out <= 32'h04000000;
             90:out <= 32'h3c000000;
             91:out <= 32'h00000000;
             92:out <= 32'h03000000;
             93:out <= 32'h15000000;
             94:out <= 32'h1b000000;
             95:out <= 32'h69666973;
             96:out <= 32'h722c6576;
             97:out <= 32'h656b636f;
             98:out <= 32'h72003074;
             99:out <= 32'h76637369;
             100:out <= 32'h00000000;
             101:out <= 32'h03000000;
             102:out <= 32'h04000000;
             103:out <= 32'h4c000000;
             104:out <= 32'h00757063;
             105:out <= 32'h03000000;
             106:out <= 32'h04000000;
             107:out <= 32'h58000000;
             108:out <= 32'h40000000;
             109:out <= 32'h03000000;
             110:out <= 32'h04000000;
             111:out <= 32'h6b000000;
             112:out <= 32'h40000000;
             113:out <= 32'h03000000;
             114:out <= 32'h04000000;
             115:out <= 32'h78000000;
             116:out <= 32'h00100000;
             117:out <= 32'h03000000;
             118:out <= 32'h04000000;
             119:out <= 32'h85000000;
             120:out <= 32'h00000000;
             121:out <= 32'h03000000;
             122:out <= 32'h09000000;
             123:out <= 32'h89000000;
             124:out <= 32'h32337672;
             125:out <= 32'h63616d69;
             126:out <= 32'h00000000;
             127:out <= 32'h03000000;
             128:out <= 32'h04000000;
             129:out <= 32'h93000000;
             130:out <= 32'h01000000;
             131:out <= 32'h03000000;
             132:out <= 32'h05000000;
             133:out <= 32'h9f000000;
             134:out <= 32'h79616b6f;
             135:out <= 32'h00000000;
             136:out <= 32'h03000000;
             137:out <= 32'h04000000;
             138:out <= 32'ha6000000;
             139:out <= 32'h00800000;
             140:out <= 32'h01000000;
             141:out <= 32'h65746e69;
             142:out <= 32'h70757272;
             143:out <= 32'h6f632d74;
             144:out <= 32'h6f72746e;
             145:out <= 32'h72656c6c;
             146:out <= 32'h00000000;
             147:out <= 32'h03000000;
             148:out <= 32'h04000000;
             149:out <= 32'hb9000000;
             150:out <= 32'h01000000;
             151:out <= 32'h03000000;
             152:out <= 32'h0f000000;
             153:out <= 32'h1b000000;
             154:out <= 32'h63736972;
             155:out <= 32'h70632c76;
             156:out <= 32'h6e692d75;
             157:out <= 32'h00006374;
             158:out <= 32'h03000000;
             159:out <= 32'h00000000;
             160:out <= 32'hca000000;
             161:out <= 32'h03000000;
             162:out <= 32'h04000000;
             163:out <= 32'hdf000000;
             164:out <= 32'h03000000;
             165:out <= 32'h03000000;
             166:out <= 32'h04000000;
             167:out <= 32'he5000000;
             168:out <= 32'h03000000;
             169:out <= 32'h02000000;
             170:out <= 32'h02000000;
             171:out <= 32'h02000000;
             172:out <= 32'h01000000;
             173:out <= 32'h00636f73;
             174:out <= 32'h03000000;
             175:out <= 32'h04000000;
             176:out <= 32'h00000000;
             177:out <= 32'h01000000;
             178:out <= 32'h03000000;
             179:out <= 32'h04000000;
             180:out <= 32'h0f000000;
             181:out <= 32'h01000000;
             182:out <= 32'h03000000;
             183:out <= 32'h2c000000;
             184:out <= 32'h1b000000;
             185:out <= 32'h65657266;
             186:out <= 32'h70696863;
             187:out <= 32'h6f722c73;
             188:out <= 32'h74656b63;
             189:out <= 32'h70696863;
             190:out <= 32'h6b6e752d;
             191:out <= 32'h6e776f6e;
             192:out <= 32'h636f732d;
             193:out <= 32'h6d697300;
             194:out <= 32'h2d656c70;
             195:out <= 32'h00737562;
             196:out <= 32'h03000000;
             197:out <= 32'h00000000;
             198:out <= 32'hed000000;
             199:out <= 32'h01000000;
             200:out <= 32'h406e6f61;
             201:out <= 32'h30303031;
             202:out <= 32'h30303030;
             203:out <= 32'h00000000;
             204:out <= 32'h03000000;
             205:out <= 32'h0c000000;
             206:out <= 32'h1b000000;
             207:out <= 32'h69666973;
             208:out <= 32'h612c6576;
             209:out <= 32'h00306e6f;
             210:out <= 32'h03000000;
             211:out <= 32'h04000000;
             212:out <= 32'hf4000000;
             213:out <= 32'h02000000;
             214:out <= 32'h03000000;
             215:out <= 32'h08000000;
             216:out <= 32'h05010000;
             217:out <= 32'h01000000;
             218:out <= 32'h02000000;
             219:out <= 32'h03000000;
             220:out <= 32'h08000000;
             221:out <= 32'h85000000;
             222:out <= 32'h00000010;
             223:out <= 32'h00100000;
             224:out <= 32'h03000000;
             225:out <= 32'h08000000;
             226:out <= 32'h10010000;
             227:out <= 32'h746e6f63;
             228:out <= 32'h006c6f72;
             229:out <= 32'h02000000;
             230:out <= 32'h01000000;
             231:out <= 32'h6e696c63;
             232:out <= 32'h30324074;
             233:out <= 32'h30303030;
             234:out <= 32'h00000030;
             235:out <= 32'h03000000;
             236:out <= 32'h0d000000;
             237:out <= 32'h1b000000;
             238:out <= 32'h63736972;
             239:out <= 32'h6c632c76;
             240:out <= 32'h30746e69;
             241:out <= 32'h00000000;
             242:out <= 32'h03000000;
             243:out <= 32'h10000000;
             244:out <= 32'h1a010000;
             245:out <= 32'h03000000;
             246:out <= 32'h03000000;
             247:out <= 32'h03000000;
             248:out <= 32'h07000000;
             249:out <= 32'h03000000;
             250:out <= 32'h08000000;
             251:out <= 32'h85000000;
             252:out <= 32'h00000002;
             253:out <= 32'h00000100;
             254:out <= 32'h03000000;
             255:out <= 32'h08000000;
             256:out <= 32'h10010000;
             257:out <= 32'h746e6f63;
             258:out <= 32'h006c6f72;
             259:out <= 32'h02000000;
             260:out <= 32'h01000000;
             261:out <= 32'h75626564;
             262:out <= 32'h6f632d67;
             263:out <= 32'h6f72746e;
             264:out <= 32'h72656c6c;
             265:out <= 32'h00003040;
             266:out <= 32'h03000000;
             267:out <= 32'h21000000;
             268:out <= 32'h1b000000;
             269:out <= 32'h69666973;
             270:out <= 32'h642c6576;
             271:out <= 32'h67756265;
             272:out <= 32'h3331302d;
             273:out <= 32'h73697200;
             274:out <= 32'h642c7663;
             275:out <= 32'h67756265;
             276:out <= 32'h3331302d;
             277:out <= 32'h00000000;
             278:out <= 32'h03000000;
             279:out <= 32'h08000000;
             280:out <= 32'h1a010000;
             281:out <= 32'h03000000;
             282:out <= 32'hffff0000;
             283:out <= 32'h03000000;
             284:out <= 32'h08000000;
             285:out <= 32'h85000000;
             286:out <= 32'h00000000;
             287:out <= 32'h00100000;
             288:out <= 32'h03000000;
             289:out <= 32'h08000000;
             290:out <= 32'h10010000;
             291:out <= 32'h746e6f63;
             292:out <= 32'h006c6f72;
             293:out <= 32'h02000000;
             294:out <= 32'h01000000;
             295:out <= 32'h6d697464;
             296:out <= 32'h30303840;
             297:out <= 32'h30303030;
             298:out <= 32'h00000030;
             299:out <= 32'h03000000;
             300:out <= 32'h0d000000;
             301:out <= 32'h1b000000;
             302:out <= 32'h69666973;
             303:out <= 32'h642c6576;
             304:out <= 32'h306d6974;
             305:out <= 32'h00000000;
             306:out <= 32'h03000000;
             307:out <= 32'h08000000;
             308:out <= 32'h85000000;
             309:out <= 32'h00000080;
             310:out <= 32'h00400000;
             311:out <= 32'h03000000;
             312:out <= 32'h04000000;
             313:out <= 32'h10010000;
             314:out <= 32'h006d656d;
             315:out <= 32'h03000000;
             316:out <= 32'h04000000;
             317:out <= 32'hdf000000;
             318:out <= 32'h01000000;
             319:out <= 32'h03000000;
             320:out <= 32'h04000000;
             321:out <= 32'he5000000;
             322:out <= 32'h01000000;
             323:out <= 32'h02000000;
             324:out <= 32'h01000000;
             325:out <= 32'h6f727265;
             326:out <= 32'h65642d72;
             327:out <= 32'h65636976;
             328:out <= 32'h30303340;
             329:out <= 32'h00000030;
             330:out <= 32'h03000000;
             331:out <= 32'h0e000000;
             332:out <= 32'h1b000000;
             333:out <= 32'h69666973;
             334:out <= 32'h652c6576;
             335:out <= 32'h726f7272;
             336:out <= 32'h00000030;
             337:out <= 32'h03000000;
             338:out <= 32'h08000000;
             339:out <= 32'h85000000;
             340:out <= 32'h00300000;
             341:out <= 32'h00100000;
             342:out <= 32'h02000000;
             343:out <= 32'h01000000;
             344:out <= 32'h6f697067;
             345:out <= 32'h30303140;
             346:out <= 32'h30303231;
             347:out <= 32'h00000030;
             348:out <= 32'h03000000;
             349:out <= 32'h04000000;
             350:out <= 32'h2e010000;
             351:out <= 32'h02000000;
             352:out <= 32'h03000000;
             353:out <= 32'h04000000;
             354:out <= 32'hb9000000;
             355:out <= 32'h02000000;
             356:out <= 32'h03000000;
             357:out <= 32'h0d000000;
             358:out <= 32'h1b000000;
             359:out <= 32'h69666973;
             360:out <= 32'h672c6576;
             361:out <= 32'h306f6970;
             362:out <= 32'h00000000;
             363:out <= 32'h03000000;
             364:out <= 32'h00000000;
             365:out <= 32'h3a010000;
             366:out <= 32'h03000000;
             367:out <= 32'h00000000;
             368:out <= 32'hca000000;
             369:out <= 32'h03000000;
             370:out <= 32'h04000000;
             371:out <= 32'hf4000000;
             372:out <= 32'h02000000;
             373:out <= 32'h03000000;
             374:out <= 32'h80000000;
             375:out <= 32'h05010000;
             376:out <= 32'h08000000;
             377:out <= 32'h09000000;
             378:out <= 32'h0a000000;
             379:out <= 32'h0b000000;
             380:out <= 32'h0c000000;
             381:out <= 32'h0d000000;
             382:out <= 32'h0e000000;
             383:out <= 32'h0f000000;
             384:out <= 32'h10000000;
             385:out <= 32'h11000000;
             386:out <= 32'h12000000;
             387:out <= 32'h13000000;
             388:out <= 32'h14000000;
             389:out <= 32'h15000000;
             390:out <= 32'h16000000;
             391:out <= 32'h17000000;
             392:out <= 32'h18000000;
             393:out <= 32'h19000000;
             394:out <= 32'h1a000000;
             395:out <= 32'h1b000000;
             396:out <= 32'h1c000000;
             397:out <= 32'h1d000000;
             398:out <= 32'h1e000000;
             399:out <= 32'h1f000000;
             400:out <= 32'h20000000;
             401:out <= 32'h21000000;
             402:out <= 32'h22000000;
             403:out <= 32'h23000000;
             404:out <= 32'h24000000;
             405:out <= 32'h25000000;
             406:out <= 32'h26000000;
             407:out <= 32'h27000000;
             408:out <= 32'h03000000;
             409:out <= 32'h08000000;
             410:out <= 32'h85000000;
             411:out <= 32'h00200110;
             412:out <= 32'h00100000;
             413:out <= 32'h03000000;
             414:out <= 32'h08000000;
             415:out <= 32'h10010000;
             416:out <= 32'h746e6f63;
             417:out <= 32'h006c6f72;
             418:out <= 32'h02000000;
             419:out <= 32'h01000000;
             420:out <= 32'h40633269;
             421:out <= 32'h31303031;
             422:out <= 32'h30303036;
             423:out <= 32'h00000000;
             424:out <= 32'h03000000;
             425:out <= 32'h0c000000;
             426:out <= 32'h1b000000;
             427:out <= 32'h69666973;
             428:out <= 32'h692c6576;
             429:out <= 32'h00306332;
             430:out <= 32'h03000000;
             431:out <= 32'h04000000;
             432:out <= 32'hf4000000;
             433:out <= 32'h02000000;
             434:out <= 32'h03000000;
             435:out <= 32'h04000000;
             436:out <= 32'h05010000;
             437:out <= 32'h34000000;
             438:out <= 32'h03000000;
             439:out <= 32'h08000000;
             440:out <= 32'h85000000;
             441:out <= 32'h00600110;
             442:out <= 32'h00100000;
             443:out <= 32'h03000000;
             444:out <= 32'h08000000;
             445:out <= 32'h10010000;
             446:out <= 32'h746e6f63;
             447:out <= 32'h006c6f72;
             448:out <= 32'h02000000;
             449:out <= 32'h01000000;
             450:out <= 32'h65746e69;
             451:out <= 32'h70757272;
             452:out <= 32'h6f632d74;
             453:out <= 32'h6f72746e;
             454:out <= 32'h72656c6c;
             455:out <= 32'h30306340;
             456:out <= 32'h30303030;
             457:out <= 32'h00000000;
             458:out <= 32'h03000000;
             459:out <= 32'h04000000;
             460:out <= 32'hb9000000;
             461:out <= 32'h01000000;
             462:out <= 32'h03000000;
             463:out <= 32'h0c000000;
             464:out <= 32'h1b000000;
             465:out <= 32'h63736972;
             466:out <= 32'h6c702c76;
             467:out <= 32'h00306369;
             468:out <= 32'h03000000;
             469:out <= 32'h00000000;
             470:out <= 32'hca000000;
             471:out <= 32'h03000000;
             472:out <= 32'h08000000;
             473:out <= 32'h1a010000;
             474:out <= 32'h03000000;
             475:out <= 32'h0b000000;
             476:out <= 32'h03000000;
             477:out <= 32'h08000000;
             478:out <= 32'h85000000;
             479:out <= 32'h0000000c;
             480:out <= 32'h00000004;
             481:out <= 32'h03000000;
             482:out <= 32'h08000000;
             483:out <= 32'h10010000;
             484:out <= 32'h746e6f63;
             485:out <= 32'h006c6f72;
             486:out <= 32'h03000000;
             487:out <= 32'h04000000;
             488:out <= 32'h4a010000;
             489:out <= 32'h07000000;
             490:out <= 32'h03000000;
             491:out <= 32'h04000000;
             492:out <= 32'h5d010000;
             493:out <= 32'h34000000;
             494:out <= 32'h03000000;
             495:out <= 32'h04000000;
             496:out <= 32'hdf000000;
             497:out <= 32'h02000000;
             498:out <= 32'h03000000;
             499:out <= 32'h04000000;
             500:out <= 32'he5000000;
             501:out <= 32'h02000000;
             502:out <= 32'h02000000;
             503:out <= 32'h01000000;
             504:out <= 32'h406d7770;
             505:out <= 32'h31303031;
             506:out <= 32'h30303035;
             507:out <= 32'h00000000;
             508:out <= 32'h03000000;
             509:out <= 32'h0c000000;
             510:out <= 32'h1b000000;
             511:out <= 32'h69666973;
             512:out <= 32'h702c6576;
             513:out <= 32'h00306d77;
             514:out <= 32'h03000000;
             515:out <= 32'h04000000;
             516:out <= 32'hf4000000;
             517:out <= 32'h02000000;
             518:out <= 32'h03000000;
             519:out <= 32'h10000000;
             520:out <= 32'h05010000;
             521:out <= 32'h28000000;
             522:out <= 32'h29000000;
             523:out <= 32'h2a000000;
             524:out <= 32'h2b000000;
             525:out <= 32'h03000000;
             526:out <= 32'h08000000;
             527:out <= 32'h85000000;
             528:out <= 32'h00500110;
             529:out <= 32'h00100000;
             530:out <= 32'h03000000;
             531:out <= 32'h08000000;
             532:out <= 32'h10010000;
             533:out <= 32'h746e6f63;
             534:out <= 32'h006c6f72;
             535:out <= 32'h02000000;
             536:out <= 32'h01000000;
             537:out <= 32'h406d7770;
             538:out <= 32'h32303031;
             539:out <= 32'h30303035;
             540:out <= 32'h00000000;
             541:out <= 32'h03000000;
             542:out <= 32'h0c000000;
             543:out <= 32'h1b000000;
             544:out <= 32'h69666973;
             545:out <= 32'h702c6576;
             546:out <= 32'h00306d77;
             547:out <= 32'h03000000;
             548:out <= 32'h04000000;
             549:out <= 32'hf4000000;
             550:out <= 32'h02000000;
             551:out <= 32'h03000000;
             552:out <= 32'h10000000;
             553:out <= 32'h05010000;
             554:out <= 32'h2c000000;
             555:out <= 32'h2d000000;
             556:out <= 32'h2e000000;
             557:out <= 32'h2f000000;
             558:out <= 32'h03000000;
             559:out <= 32'h08000000;
             560:out <= 32'h85000000;
             561:out <= 32'h00500210;
             562:out <= 32'h00100000;
             563:out <= 32'h03000000;
             564:out <= 32'h08000000;
             565:out <= 32'h10010000;
             566:out <= 32'h746e6f63;
             567:out <= 32'h006c6f72;
             568:out <= 32'h02000000;
             569:out <= 32'h01000000;
             570:out <= 32'h406d7770;
             571:out <= 32'h33303031;
             572:out <= 32'h30303035;
             573:out <= 32'h00000000;
             574:out <= 32'h03000000;
             575:out <= 32'h0c000000;
             576:out <= 32'h1b000000;
             577:out <= 32'h69666973;
             578:out <= 32'h702c6576;
             579:out <= 32'h00306d77;
             580:out <= 32'h03000000;
             581:out <= 32'h04000000;
             582:out <= 32'hf4000000;
             583:out <= 32'h02000000;
             584:out <= 32'h03000000;
             585:out <= 32'h10000000;
             586:out <= 32'h05010000;
             587:out <= 32'h30000000;
             588:out <= 32'h31000000;
             589:out <= 32'h32000000;
             590:out <= 32'h33000000;
             591:out <= 32'h03000000;
             592:out <= 32'h08000000;
             593:out <= 32'h85000000;
             594:out <= 32'h00500310;
             595:out <= 32'h00100000;
             596:out <= 32'h03000000;
             597:out <= 32'h08000000;
             598:out <= 32'h10010000;
             599:out <= 32'h746e6f63;
             600:out <= 32'h006c6f72;
             601:out <= 32'h02000000;
             602:out <= 32'h01000000;
             603:out <= 32'h406d6f72;
             604:out <= 32'h30303031;
             605:out <= 32'h00000030;
             606:out <= 32'h03000000;
             607:out <= 32'h10000000;
             608:out <= 32'h1b000000;
             609:out <= 32'h69666973;
             610:out <= 32'h6d2c6576;
             611:out <= 32'h726b7361;
             612:out <= 32'h00306d6f;
             613:out <= 32'h03000000;
             614:out <= 32'h08000000;
             615:out <= 32'h85000000;
             616:out <= 32'h00000100;
             617:out <= 32'h00200000;
             618:out <= 32'h03000000;
             619:out <= 32'h04000000;
             620:out <= 32'h10010000;
             621:out <= 32'h006d656d;
             622:out <= 32'h02000000;
             623:out <= 32'h01000000;
             624:out <= 32'h69726573;
             625:out <= 32'h31406c61;
             626:out <= 32'h33313030;
             627:out <= 32'h00303030;
             628:out <= 32'h03000000;
             629:out <= 32'h0d000000;
             630:out <= 32'h1b000000;
             631:out <= 32'h69666973;
             632:out <= 32'h752c6576;
             633:out <= 32'h30747261;
             634:out <= 32'h00000000;
             635:out <= 32'h03000000;
             636:out <= 32'h04000000;
             637:out <= 32'hf4000000;
             638:out <= 32'h02000000;
             639:out <= 32'h03000000;
             640:out <= 32'h04000000;
             641:out <= 32'h05010000;
             642:out <= 32'h03000000;
             643:out <= 32'h03000000;
             644:out <= 32'h08000000;
             645:out <= 32'h85000000;
             646:out <= 32'h00300110;
             647:out <= 32'h00100000;
             648:out <= 32'h03000000;
             649:out <= 32'h08000000;
             650:out <= 32'h10010000;
             651:out <= 32'h746e6f63;
             652:out <= 32'h006c6f72;
             653:out <= 32'h02000000;
             654:out <= 32'h01000000;
             655:out <= 32'h69726573;
             656:out <= 32'h31406c61;
             657:out <= 32'h33323030;
             658:out <= 32'h00303030;
             659:out <= 32'h03000000;
             660:out <= 32'h0d000000;
             661:out <= 32'h1b000000;
             662:out <= 32'h69666973;
             663:out <= 32'h752c6576;
             664:out <= 32'h30747261;
             665:out <= 32'h00000000;
             666:out <= 32'h03000000;
             667:out <= 32'h04000000;
             668:out <= 32'hf4000000;
             669:out <= 32'h02000000;
             670:out <= 32'h03000000;
             671:out <= 32'h04000000;
             672:out <= 32'h05010000;
             673:out <= 32'h04000000;
             674:out <= 32'h03000000;
             675:out <= 32'h08000000;
             676:out <= 32'h85000000;
             677:out <= 32'h00300210;
             678:out <= 32'h00100000;
             679:out <= 32'h03000000;
             680:out <= 32'h08000000;
             681:out <= 32'h10010000;
             682:out <= 32'h746e6f63;
             683:out <= 32'h006c6f72;
             684:out <= 32'h02000000;
             685:out <= 32'h01000000;
             686:out <= 32'h40697073;
             687:out <= 32'h31303031;
             688:out <= 32'h30303034;
             689:out <= 32'h00000000;
             690:out <= 32'h03000000;
             691:out <= 32'h04000000;
             692:out <= 32'h00000000;
             693:out <= 32'h01000000;
             694:out <= 32'h03000000;
             695:out <= 32'h04000000;
             696:out <= 32'h0f000000;
             697:out <= 32'h00000000;
             698:out <= 32'h03000000;
             699:out <= 32'h0c000000;
             700:out <= 32'h1b000000;
             701:out <= 32'h69666973;
             702:out <= 32'h732c6576;
             703:out <= 32'h00306970;
             704:out <= 32'h03000000;
             705:out <= 32'h04000000;
             706:out <= 32'hf4000000;
             707:out <= 32'h02000000;
             708:out <= 32'h03000000;
             709:out <= 32'h04000000;
             710:out <= 32'h05010000;
             711:out <= 32'h05000000;
             712:out <= 32'h03000000;
             713:out <= 32'h10000000;
             714:out <= 32'h85000000;
             715:out <= 32'h00400110;
             716:out <= 32'h00100000;
             717:out <= 32'h00000020;
             718:out <= 32'h00000020;
             719:out <= 32'h03000000;
             720:out <= 32'h0c000000;
             721:out <= 32'h10010000;
             722:out <= 32'h746e6f63;
             723:out <= 32'h006c6f72;
             724:out <= 32'h006d656d;
             725:out <= 32'h02000000;
             726:out <= 32'h01000000;
             727:out <= 32'h40697073;
             728:out <= 32'h32303031;
             729:out <= 32'h30303034;
             730:out <= 32'h00000000;
             731:out <= 32'h03000000;
             732:out <= 32'h04000000;
             733:out <= 32'h00000000;
             734:out <= 32'h01000000;
             735:out <= 32'h03000000;
             736:out <= 32'h04000000;
             737:out <= 32'h0f000000;
             738:out <= 32'h00000000;
             739:out <= 32'h03000000;
             740:out <= 32'h0c000000;
             741:out <= 32'h1b000000;
             742:out <= 32'h69666973;
             743:out <= 32'h732c6576;
             744:out <= 32'h00306970;
             745:out <= 32'h03000000;
             746:out <= 32'h04000000;
             747:out <= 32'hf4000000;
             748:out <= 32'h02000000;
             749:out <= 32'h03000000;
             750:out <= 32'h04000000;
             751:out <= 32'h05010000;
             752:out <= 32'h06000000;
             753:out <= 32'h03000000;
             754:out <= 32'h08000000;
             755:out <= 32'h85000000;
             756:out <= 32'h00400210;
             757:out <= 32'h00100000;
             758:out <= 32'h03000000;
             759:out <= 32'h08000000;
             760:out <= 32'h10010000;
             761:out <= 32'h746e6f63;
             762:out <= 32'h006c6f72;
             763:out <= 32'h02000000;
             764:out <= 32'h01000000;
             765:out <= 32'h40697073;
             766:out <= 32'h33303031;
             767:out <= 32'h30303034;
             768:out <= 32'h00000000;
             769:out <= 32'h03000000;
             770:out <= 32'h04000000;
             771:out <= 32'h00000000;
             772:out <= 32'h01000000;
             773:out <= 32'h03000000;
             774:out <= 32'h04000000;
             775:out <= 32'h0f000000;
             776:out <= 32'h00000000;
             777:out <= 32'h03000000;
             778:out <= 32'h0c000000;
             779:out <= 32'h1b000000;
             780:out <= 32'h69666973;
             781:out <= 32'h732c6576;
             782:out <= 32'h00306970;
             783:out <= 32'h03000000;
             784:out <= 32'h04000000;
             785:out <= 32'hf4000000;
             786:out <= 32'h02000000;
             787:out <= 32'h03000000;
             788:out <= 32'h04000000;
             789:out <= 32'h05010000;
             790:out <= 32'h07000000;
             791:out <= 32'h03000000;
             792:out <= 32'h08000000;
             793:out <= 32'h85000000;
             794:out <= 32'h00400310;
             795:out <= 32'h00100000;
             796:out <= 32'h03000000;
             797:out <= 32'h08000000;
             798:out <= 32'h10010000;
             799:out <= 32'h746e6f63;
             800:out <= 32'h006c6f72;
             801:out <= 32'h02000000;
             802:out <= 32'h02000000;
             803:out <= 32'h02000000;
             804:out <= 32'h09000000;
             805:out <= 32'h64646123;
             806:out <= 32'h73736572;
             807:out <= 32'h6c65632d;
             808:out <= 32'h2300736c;
             809:out <= 32'h657a6973;
             810:out <= 32'h6c65632d;
             811:out <= 32'h6300736c;
             812:out <= 32'h61706d6f;
             813:out <= 32'h6c626974;
             814:out <= 32'h6f6d0065;
             815:out <= 32'h006c6564;
             816:out <= 32'h69726573;
             817:out <= 32'h00306c61;
             818:out <= 32'h69726573;
             819:out <= 32'h00316c61;
             820:out <= 32'h636f6c63;
             821:out <= 32'h72662d6b;
             822:out <= 32'h65757165;
             823:out <= 32'h0079636e;
             824:out <= 32'h69766564;
             825:out <= 32'h745f6563;
             826:out <= 32'h00657079;
             827:out <= 32'h61632d69;
             828:out <= 32'h2d656863;
             829:out <= 32'h636f6c62;
             830:out <= 32'h69732d6b;
             831:out <= 32'h6900657a;
             832:out <= 32'h6361632d;
             833:out <= 32'h732d6568;
             834:out <= 32'h00737465;
             835:out <= 32'h61632d69;
             836:out <= 32'h2d656863;
             837:out <= 32'h657a6973;
             838:out <= 32'h67657200;
             839:out <= 32'h73697200;
             840:out <= 32'h692c7663;
             841:out <= 32'h73006173;
             842:out <= 32'h76696669;
             843:out <= 32'h74642c65;
             844:out <= 32'h73006d69;
             845:out <= 32'h75746174;
             846:out <= 32'h69740073;
             847:out <= 32'h6162656d;
             848:out <= 32'h662d6573;
             849:out <= 32'h75716572;
             850:out <= 32'h79636e65;
             851:out <= 32'h6e692300;
             852:out <= 32'h72726574;
             853:out <= 32'h2d747075;
             854:out <= 32'h6c6c6563;
             855:out <= 32'h6e690073;
             856:out <= 32'h72726574;
             857:out <= 32'h2d747075;
             858:out <= 32'h746e6f63;
             859:out <= 32'h6c6c6f72;
             860:out <= 32'h6c007265;
             861:out <= 32'h78756e69;
             862:out <= 32'h6168702c;
             863:out <= 32'h656c646e;
             864:out <= 32'h6e617200;
             865:out <= 32'h00736567;
             866:out <= 32'h65746e69;
             867:out <= 32'h70757272;
             868:out <= 32'h61702d74;
             869:out <= 32'h746e6572;
             870:out <= 32'h746e6900;
             871:out <= 32'h75727265;
             872:out <= 32'h00737470;
             873:out <= 32'h2d676572;
             874:out <= 32'h656d616e;
             875:out <= 32'h6e690073;
             876:out <= 32'h72726574;
             877:out <= 32'h73747075;
             878:out <= 32'h7478652d;
             879:out <= 32'h65646e65;
             880:out <= 32'h67230064;
             881:out <= 32'h2d6f6970;
             882:out <= 32'h6c6c6563;
             883:out <= 32'h70670073;
             884:out <= 32'h632d6f69;
             885:out <= 32'h72746e6f;
             886:out <= 32'h656c6c6f;
             887:out <= 32'h69720072;
             888:out <= 32'h2c766373;
             889:out <= 32'h2d78616d;
             890:out <= 32'h6f697270;
             891:out <= 32'h79746972;
             892:out <= 32'h73697200;
             893:out <= 32'h6e2c7663;
             894:out <= 32'h00766564;
             895:out <= 32'h00000000;
             896:out <= 32'h00000000;
             897:out <= 32'h00000000;
             898:out <= 32'h00000000;
             899:out <= 32'h00000000;
             900:out <= 32'h00000000;
             901:out <= 32'h00000000;
             902:out <= 32'h00000000;
             903:out <= 32'h00000000;
             904:out <= 32'h00000000;
             905:out <= 32'h00000000;
             906:out <= 32'h00000000;
             907:out <= 32'h00000000;
             908:out <= 32'h00000000;
             909:out <= 32'h00000000;
             910:out <= 32'h00000000;
             911:out <= 32'h00000000;
             912:out <= 32'h00000000;
             913:out <= 32'h00000000;
             914:out <= 32'h00000000;
             915:out <= 32'h00000000;
             916:out <= 32'h00000000;
             917:out <= 32'h00000000;
             918:out <= 32'h00000000;
             919:out <= 32'h00000000;
             920:out <= 32'h00000000;
             921:out <= 32'h00000000;
             922:out <= 32'h00000000;
             923:out <= 32'h00000000;
             924:out <= 32'h00000000;
             925:out <= 32'h00000000;
             926:out <= 32'h00000000;
             927:out <= 32'h00000000;
             928:out <= 32'h00000000;
             929:out <= 32'h00000000;
             930:out <= 32'h00000000;
             931:out <= 32'h00000000;
             932:out <= 32'h00000000;
             933:out <= 32'h00000000;
             934:out <= 32'h00000000;
             935:out <= 32'h00000000;
             936:out <= 32'h00000000;
             937:out <= 32'h00000000;
             938:out <= 32'h00000000;
             939:out <= 32'h00000000;
             940:out <= 32'h00000000;
             941:out <= 32'h00000000;
             942:out <= 32'h00000000;
             943:out <= 32'h00000000;
             944:out <= 32'h00000000;
             945:out <= 32'h00000000;
             946:out <= 32'h00000000;
             947:out <= 32'h00000000;
             948:out <= 32'h00000000;
             949:out <= 32'h00000000;
             950:out <= 32'h00000000;
             951:out <= 32'h00000000;
             952:out <= 32'h00000000;
             953:out <= 32'h00000000;
             954:out <= 32'h00000000;
             955:out <= 32'h00000000;
             956:out <= 32'h00000000;
             957:out <= 32'h00000000;
             958:out <= 32'h00000000;
             959:out <= 32'h00000000;
             960:out <= 32'h00000000;
             961:out <= 32'h00000000;
             962:out <= 32'h00000000;
             963:out <= 32'h00000000;
             964:out <= 32'h00000000;
             965:out <= 32'h00000000;
             966:out <= 32'h00000000;
             967:out <= 32'h00000000;
             968:out <= 32'h00000000;
             969:out <= 32'h00000000;
             970:out <= 32'h00000000;
             971:out <= 32'h00000000;
             972:out <= 32'h00000000;
             973:out <= 32'h00000000;
             974:out <= 32'h00000000;
             975:out <= 32'h00000000;
             976:out <= 32'h00000000;
             977:out <= 32'h00000000;
             978:out <= 32'h00000000;
             979:out <= 32'h00000000;
             980:out <= 32'h00000000;
             981:out <= 32'h00000000;
             982:out <= 32'h00000000;
             983:out <= 32'h00000000;
             984:out <= 32'h00000000;
             985:out <= 32'h00000000;
             986:out <= 32'h00000000;
             987:out <= 32'h00000000;
             988:out <= 32'h00000000;
             989:out <= 32'h00000000;
             990:out <= 32'h00000000;
             991:out <= 32'h00000000;
             992:out <= 32'h00000000;
             993:out <= 32'h00000000;
             994:out <= 32'h00000000;
             995:out <= 32'h00000000;
             996:out <= 32'h00000000;
             997:out <= 32'h00000000;
             998:out <= 32'h00000000;
             999:out <= 32'h00000000;
             1000:out <= 32'h00000000;
             1001:out <= 32'h00000000;
             1002:out <= 32'h00000000;
             1003:out <= 32'h00000000;
             1004:out <= 32'h00000000;
             1005:out <= 32'h00000000;
             1006:out <= 32'h00000000;
             1007:out <= 32'h00000000;
             1008:out <= 32'h00000000;
             1009:out <= 32'h00000000;
             1010:out <= 32'h00000000;
             1011:out <= 32'h00000000;
             1012:out <= 32'h00000000;
             1013:out <= 32'h00000000;
             1014:out <= 32'h00000000;
             1015:out <= 32'h00000000;
             1016:out <= 32'h00000000;
             1017:out <= 32'h00000000;
             1018:out <= 32'h00000000;
             1019:out <= 32'h00000000;
             1020:out <= 32'h00000000;
             1021:out <= 32'h00000000;
             1022:out <= 32'h00000000;
             1023:out <= 32'h00000000;
             1024:out <= 32'h00000000;
             1025:out <= 32'h00000000;
             1026:out <= 32'h00000000;
             1027:out <= 32'h00000000;
             1028:out <= 32'h00000000;
             1029:out <= 32'h00000000;
             1030:out <= 32'h00000000;
             1031:out <= 32'h00000000;
             1032:out <= 32'h00000000;
             1033:out <= 32'h00000000;
             1034:out <= 32'h00000000;
             1035:out <= 32'h00000000;
             1036:out <= 32'h00000000;
             1037:out <= 32'h00000000;
             1038:out <= 32'h00000000;
             1039:out <= 32'h00000000;
             1040:out <= 32'h00000000;
             1041:out <= 32'h00000000;
             1042:out <= 32'h00000000;
             1043:out <= 32'h00000000;
             1044:out <= 32'h00000000;
             1045:out <= 32'h00000000;
             1046:out <= 32'h00000000;
             1047:out <= 32'h00000000;
             1048:out <= 32'h00000000;
             1049:out <= 32'h00000000;
             1050:out <= 32'h00000000;
             1051:out <= 32'h00000000;
             1052:out <= 32'h00000000;
             1053:out <= 32'h00000000;
             1054:out <= 32'h00000000;
             1055:out <= 32'h00000000;
             1056:out <= 32'h00000000;
             1057:out <= 32'h00000000;
             1058:out <= 32'h00000000;
             1059:out <= 32'h00000000;
             1060:out <= 32'h00000000;
             1061:out <= 32'h00000000;
             1062:out <= 32'h00000000;
             1063:out <= 32'h00000000;
             1064:out <= 32'h00000000;
             1065:out <= 32'h00000000;
             1066:out <= 32'h00000000;
             1067:out <= 32'h00000000;
             1068:out <= 32'h00000000;
             1069:out <= 32'h00000000;
             1070:out <= 32'h00000000;
             1071:out <= 32'h00000000;
             1072:out <= 32'h00000000;
             1073:out <= 32'h00000000;
             1074:out <= 32'h00000000;
             1075:out <= 32'h00000000;
             1076:out <= 32'h00000000;
             1077:out <= 32'h00000000;
             1078:out <= 32'h00000000;
             1079:out <= 32'h00000000;
             1080:out <= 32'h00000000;
             1081:out <= 32'h00000000;
             1082:out <= 32'h00000000;
             1083:out <= 32'h00000000;
             1084:out <= 32'h00000000;
             1085:out <= 32'h00000000;
             1086:out <= 32'h00000000;
             1087:out <= 32'h00000000;
             1088:out <= 32'h00000000;
             1089:out <= 32'h00000000;
             1090:out <= 32'h00000000;
             1091:out <= 32'h00000000;
             1092:out <= 32'h00000000;
             1093:out <= 32'h00000000;
             1094:out <= 32'h00000000;
             1095:out <= 32'h00000000;
             1096:out <= 32'h00000000;
             1097:out <= 32'h00000000;
             1098:out <= 32'h00000000;
             1099:out <= 32'h00000000;
             1100:out <= 32'h00000000;
             1101:out <= 32'h00000000;
             1102:out <= 32'h00000000;
             1103:out <= 32'h00000000;
             1104:out <= 32'h00000000;
             1105:out <= 32'h00000000;
             1106:out <= 32'h00000000;
             1107:out <= 32'h00000000;
             1108:out <= 32'h00000000;
             1109:out <= 32'h00000000;
             1110:out <= 32'h00000000;
             1111:out <= 32'h00000000;
             1112:out <= 32'h00000000;
             1113:out <= 32'h00000000;
             1114:out <= 32'h00000000;
             1115:out <= 32'h00000000;
             1116:out <= 32'h00000000;
             1117:out <= 32'h00000000;
             1118:out <= 32'h00000000;
             1119:out <= 32'h00000000;
             1120:out <= 32'h00000000;
             1121:out <= 32'h00000000;
             1122:out <= 32'h00000000;
             1123:out <= 32'h00000000;
             1124:out <= 32'h00000000;
             1125:out <= 32'h00000000;
             1126:out <= 32'h00000000;
             1127:out <= 32'h00000000;
             1128:out <= 32'h00000000;
             1129:out <= 32'h00000000;
             1130:out <= 32'h00000000;
             1131:out <= 32'h00000000;
             1132:out <= 32'h00000000;
             1133:out <= 32'h00000000;
             1134:out <= 32'h00000000;
             1135:out <= 32'h00000000;
             1136:out <= 32'h00000000;
             1137:out <= 32'h00000000;
             1138:out <= 32'h00000000;
             1139:out <= 32'h00000000;
             1140:out <= 32'h00000000;
             1141:out <= 32'h00000000;
             1142:out <= 32'h00000000;
             1143:out <= 32'h00000000;
             1144:out <= 32'h00000000;
             1145:out <= 32'h00000000;
             1146:out <= 32'h00000000;
             1147:out <= 32'h00000000;
             1148:out <= 32'h00000000;
             1149:out <= 32'h00000000;
             1150:out <= 32'h00000000;
             1151:out <= 32'h00000000;
             1152:out <= 32'h00000000;
             1153:out <= 32'h00000000;
             1154:out <= 32'h00000000;
             1155:out <= 32'h00000000;
             1156:out <= 32'h00000000;
             1157:out <= 32'h00000000;
             1158:out <= 32'h00000000;
             1159:out <= 32'h00000000;
             1160:out <= 32'h00000000;
             1161:out <= 32'h00000000;
             1162:out <= 32'h00000000;
             1163:out <= 32'h00000000;
             1164:out <= 32'h00000000;
             1165:out <= 32'h00000000;
             1166:out <= 32'h00000000;
             1167:out <= 32'h00000000;
             1168:out <= 32'h00000000;
             1169:out <= 32'h00000000;
             1170:out <= 32'h00000000;
             1171:out <= 32'h00000000;
             1172:out <= 32'h00000000;
             1173:out <= 32'h00000000;
             1174:out <= 32'h00000000;
             1175:out <= 32'h00000000;
             1176:out <= 32'h00000000;
             1177:out <= 32'h00000000;
             1178:out <= 32'h00000000;
             1179:out <= 32'h00000000;
             1180:out <= 32'h00000000;
             1181:out <= 32'h00000000;
             1182:out <= 32'h00000000;
             1183:out <= 32'h00000000;
             1184:out <= 32'h00000000;
             1185:out <= 32'h00000000;
             1186:out <= 32'h00000000;
             1187:out <= 32'h00000000;
             1188:out <= 32'h00000000;
             1189:out <= 32'h00000000;
             1190:out <= 32'h00000000;
             1191:out <= 32'h00000000;
             1192:out <= 32'h00000000;
             1193:out <= 32'h00000000;
             1194:out <= 32'h00000000;
             1195:out <= 32'h00000000;
             1196:out <= 32'h00000000;
             1197:out <= 32'h00000000;
             1198:out <= 32'h00000000;
             1199:out <= 32'h00000000;
             1200:out <= 32'h00000000;
             1201:out <= 32'h00000000;
             1202:out <= 32'h00000000;
             1203:out <= 32'h00000000;
             1204:out <= 32'h00000000;
             1205:out <= 32'h00000000;
             1206:out <= 32'h00000000;
             1207:out <= 32'h00000000;
             1208:out <= 32'h00000000;
             1209:out <= 32'h00000000;
             1210:out <= 32'h00000000;
             1211:out <= 32'h00000000;
             1212:out <= 32'h00000000;
             1213:out <= 32'h00000000;
             1214:out <= 32'h00000000;
             1215:out <= 32'h00000000;
             1216:out <= 32'h00000000;
             1217:out <= 32'h00000000;
             1218:out <= 32'h00000000;
             1219:out <= 32'h00000000;
             1220:out <= 32'h00000000;
             1221:out <= 32'h00000000;
             1222:out <= 32'h00000000;
             1223:out <= 32'h00000000;
             1224:out <= 32'h00000000;
             1225:out <= 32'h00000000;
             1226:out <= 32'h00000000;
             1227:out <= 32'h00000000;
             1228:out <= 32'h00000000;
             1229:out <= 32'h00000000;
             1230:out <= 32'h00000000;
             1231:out <= 32'h00000000;
             1232:out <= 32'h00000000;
             1233:out <= 32'h00000000;
             1234:out <= 32'h00000000;
             1235:out <= 32'h00000000;
             1236:out <= 32'h00000000;
             1237:out <= 32'h00000000;
             1238:out <= 32'h00000000;
             1239:out <= 32'h00000000;
             1240:out <= 32'h00000000;
             1241:out <= 32'h00000000;
             1242:out <= 32'h00000000;
             1243:out <= 32'h00000000;
             1244:out <= 32'h00000000;
             1245:out <= 32'h00000000;
             1246:out <= 32'h00000000;
             1247:out <= 32'h00000000;
             1248:out <= 32'h00000000;
             1249:out <= 32'h00000000;
             1250:out <= 32'h00000000;
             1251:out <= 32'h00000000;
             1252:out <= 32'h00000000;
             1253:out <= 32'h00000000;
             1254:out <= 32'h00000000;
             1255:out <= 32'h00000000;
             1256:out <= 32'h00000000;
             1257:out <= 32'h00000000;
             1258:out <= 32'h00000000;
             1259:out <= 32'h00000000;
             1260:out <= 32'h00000000;
             1261:out <= 32'h00000000;
             1262:out <= 32'h00000000;
             1263:out <= 32'h00000000;
             1264:out <= 32'h00000000;
             1265:out <= 32'h00000000;
             1266:out <= 32'h00000000;
             1267:out <= 32'h00000000;
             1268:out <= 32'h00000000;
             1269:out <= 32'h00000000;
             1270:out <= 32'h00000000;
             1271:out <= 32'h00000000;
             1272:out <= 32'h00000000;
             1273:out <= 32'h00000000;
             1274:out <= 32'h00000000;
             1275:out <= 32'h00000000;
             1276:out <= 32'h00000000;
             1277:out <= 32'h00000000;
             1278:out <= 32'h00000000;
             1279:out <= 32'h00000000;
             1280:out <= 32'h00000000;
             1281:out <= 32'h00000000;
             1282:out <= 32'h00000000;
             1283:out <= 32'h00000000;
             1284:out <= 32'h00000000;
             1285:out <= 32'h00000000;
             1286:out <= 32'h00000000;
             1287:out <= 32'h00000000;
             1288:out <= 32'h00000000;
             1289:out <= 32'h00000000;
             1290:out <= 32'h00000000;
             1291:out <= 32'h00000000;
             1292:out <= 32'h00000000;
             1293:out <= 32'h00000000;
             1294:out <= 32'h00000000;
             1295:out <= 32'h00000000;
             1296:out <= 32'h00000000;
             1297:out <= 32'h00000000;
             1298:out <= 32'h00000000;
             1299:out <= 32'h00000000;
             1300:out <= 32'h00000000;
             1301:out <= 32'h00000000;
             1302:out <= 32'h00000000;
             1303:out <= 32'h00000000;
             1304:out <= 32'h00000000;
             1305:out <= 32'h00000000;
             1306:out <= 32'h00000000;
             1307:out <= 32'h00000000;
             1308:out <= 32'h00000000;
             1309:out <= 32'h00000000;
             1310:out <= 32'h00000000;
             1311:out <= 32'h00000000;
             1312:out <= 32'h00000000;
             1313:out <= 32'h00000000;
             1314:out <= 32'h00000000;
             1315:out <= 32'h00000000;
             1316:out <= 32'h00000000;
             1317:out <= 32'h00000000;
             1318:out <= 32'h00000000;
             1319:out <= 32'h00000000;
             1320:out <= 32'h00000000;
             1321:out <= 32'h00000000;
             1322:out <= 32'h00000000;
             1323:out <= 32'h00000000;
             1324:out <= 32'h00000000;
             1325:out <= 32'h00000000;
             1326:out <= 32'h00000000;
             1327:out <= 32'h00000000;
             1328:out <= 32'h00000000;
             1329:out <= 32'h00000000;
             1330:out <= 32'h00000000;
             1331:out <= 32'h00000000;
             1332:out <= 32'h00000000;
             1333:out <= 32'h00000000;
             1334:out <= 32'h00000000;
             1335:out <= 32'h00000000;
             1336:out <= 32'h00000000;
             1337:out <= 32'h00000000;
             1338:out <= 32'h00000000;
             1339:out <= 32'h00000000;
             1340:out <= 32'h00000000;
             1341:out <= 32'h00000000;
             1342:out <= 32'h00000000;
             1343:out <= 32'h00000000;
             1344:out <= 32'h00000000;
             1345:out <= 32'h00000000;
             1346:out <= 32'h00000000;
             1347:out <= 32'h00000000;
             1348:out <= 32'h00000000;
             1349:out <= 32'h00000000;
             1350:out <= 32'h00000000;
             1351:out <= 32'h00000000;
             1352:out <= 32'h00000000;
             1353:out <= 32'h00000000;
             1354:out <= 32'h00000000;
             1355:out <= 32'h00000000;
             1356:out <= 32'h00000000;
             1357:out <= 32'h00000000;
             1358:out <= 32'h00000000;
             1359:out <= 32'h00000000;
             1360:out <= 32'h00000000;
             1361:out <= 32'h00000000;
             1362:out <= 32'h00000000;
             1363:out <= 32'h00000000;
             1364:out <= 32'h00000000;
             1365:out <= 32'h00000000;
             1366:out <= 32'h00000000;
             1367:out <= 32'h00000000;
             1368:out <= 32'h00000000;
             1369:out <= 32'h00000000;
             1370:out <= 32'h00000000;
             1371:out <= 32'h00000000;
             1372:out <= 32'h00000000;
             1373:out <= 32'h00000000;
             1374:out <= 32'h00000000;
             1375:out <= 32'h00000000;
             1376:out <= 32'h00000000;
             1377:out <= 32'h00000000;
             1378:out <= 32'h00000000;
             1379:out <= 32'h00000000;
             1380:out <= 32'h00000000;
             1381:out <= 32'h00000000;
             1382:out <= 32'h00000000;
             1383:out <= 32'h00000000;
             1384:out <= 32'h00000000;
             1385:out <= 32'h00000000;
             1386:out <= 32'h00000000;
             1387:out <= 32'h00000000;
             1388:out <= 32'h00000000;
             1389:out <= 32'h00000000;
             1390:out <= 32'h00000000;
             1391:out <= 32'h00000000;
             1392:out <= 32'h00000000;
             1393:out <= 32'h00000000;
             1394:out <= 32'h00000000;
             1395:out <= 32'h00000000;
             1396:out <= 32'h00000000;
             1397:out <= 32'h00000000;
             1398:out <= 32'h00000000;
             1399:out <= 32'h00000000;
             1400:out <= 32'h00000000;
             1401:out <= 32'h00000000;
             1402:out <= 32'h00000000;
             1403:out <= 32'h00000000;
             1404:out <= 32'h00000000;
             1405:out <= 32'h00000000;
             1406:out <= 32'h00000000;
             1407:out <= 32'h00000000;
             1408:out <= 32'h00000000;
             1409:out <= 32'h00000000;
             1410:out <= 32'h00000000;
             1411:out <= 32'h00000000;
             1412:out <= 32'h00000000;
             1413:out <= 32'h00000000;
             1414:out <= 32'h00000000;
             1415:out <= 32'h00000000;
             1416:out <= 32'h00000000;
             1417:out <= 32'h00000000;
             1418:out <= 32'h00000000;
             1419:out <= 32'h00000000;
             1420:out <= 32'h00000000;
             1421:out <= 32'h00000000;
             1422:out <= 32'h00000000;
             1423:out <= 32'h00000000;
             1424:out <= 32'h00000000;
             1425:out <= 32'h00000000;
             1426:out <= 32'h00000000;
             1427:out <= 32'h00000000;
             1428:out <= 32'h00000000;
             1429:out <= 32'h00000000;
             1430:out <= 32'h00000000;
             1431:out <= 32'h00000000;
             1432:out <= 32'h00000000;
             1433:out <= 32'h00000000;
             1434:out <= 32'h00000000;
             1435:out <= 32'h00000000;
             1436:out <= 32'h00000000;
             1437:out <= 32'h00000000;
             1438:out <= 32'h00000000;
             1439:out <= 32'h00000000;
             1440:out <= 32'h00000000;
             1441:out <= 32'h00000000;
             1442:out <= 32'h00000000;
             1443:out <= 32'h00000000;
             1444:out <= 32'h00000000;
             1445:out <= 32'h00000000;
             1446:out <= 32'h00000000;
             1447:out <= 32'h00000000;
             1448:out <= 32'h00000000;
             1449:out <= 32'h00000000;
             1450:out <= 32'h00000000;
             1451:out <= 32'h00000000;
             1452:out <= 32'h00000000;
             1453:out <= 32'h00000000;
             1454:out <= 32'h00000000;
             1455:out <= 32'h00000000;
             1456:out <= 32'h00000000;
             1457:out <= 32'h00000000;
             1458:out <= 32'h00000000;
             1459:out <= 32'h00000000;
             1460:out <= 32'h00000000;
             1461:out <= 32'h00000000;
             1462:out <= 32'h00000000;
             1463:out <= 32'h00000000;
             1464:out <= 32'h00000000;
             1465:out <= 32'h00000000;
             1466:out <= 32'h00000000;
             1467:out <= 32'h00000000;
             1468:out <= 32'h00000000;
             1469:out <= 32'h00000000;
             1470:out <= 32'h00000000;
             1471:out <= 32'h00000000;
             1472:out <= 32'h00000000;
             1473:out <= 32'h00000000;
             1474:out <= 32'h00000000;
             1475:out <= 32'h00000000;
             1476:out <= 32'h00000000;
             1477:out <= 32'h00000000;
             1478:out <= 32'h00000000;
             1479:out <= 32'h00000000;
             1480:out <= 32'h00000000;
             1481:out <= 32'h00000000;
             1482:out <= 32'h00000000;
             1483:out <= 32'h00000000;
             1484:out <= 32'h00000000;
             1485:out <= 32'h00000000;
             1486:out <= 32'h00000000;
             1487:out <= 32'h00000000;
             1488:out <= 32'h00000000;
             1489:out <= 32'h00000000;
             1490:out <= 32'h00000000;
             1491:out <= 32'h00000000;
             1492:out <= 32'h00000000;
             1493:out <= 32'h00000000;
             1494:out <= 32'h00000000;
             1495:out <= 32'h00000000;
             1496:out <= 32'h00000000;
             1497:out <= 32'h00000000;
             1498:out <= 32'h00000000;
             1499:out <= 32'h00000000;
             1500:out <= 32'h00000000;
             1501:out <= 32'h00000000;
             1502:out <= 32'h00000000;
             1503:out <= 32'h00000000;
             1504:out <= 32'h00000000;
             1505:out <= 32'h00000000;
             1506:out <= 32'h00000000;
             1507:out <= 32'h00000000;
             1508:out <= 32'h00000000;
             1509:out <= 32'h00000000;
             1510:out <= 32'h00000000;
             1511:out <= 32'h00000000;
             1512:out <= 32'h00000000;
             1513:out <= 32'h00000000;
             1514:out <= 32'h00000000;
             1515:out <= 32'h00000000;
             1516:out <= 32'h00000000;
             1517:out <= 32'h00000000;
             1518:out <= 32'h00000000;
             1519:out <= 32'h00000000;
             1520:out <= 32'h00000000;
             1521:out <= 32'h00000000;
             1522:out <= 32'h00000000;
             1523:out <= 32'h00000000;
             1524:out <= 32'h00000000;
             1525:out <= 32'h00000000;
             1526:out <= 32'h00000000;
             1527:out <= 32'h00000000;
             1528:out <= 32'h00000000;
             1529:out <= 32'h00000000;
             1530:out <= 32'h00000000;
             1531:out <= 32'h00000000;
             1532:out <= 32'h00000000;
             1533:out <= 32'h00000000;
             1534:out <= 32'h00000000;
             1535:out <= 32'h00000000;
             1536:out <= 32'h00000000;
             1537:out <= 32'h00000000;
             1538:out <= 32'h00000000;
             1539:out <= 32'h00000000;
             1540:out <= 32'h00000000;
             1541:out <= 32'h00000000;
             1542:out <= 32'h00000000;
             1543:out <= 32'h00000000;
             1544:out <= 32'h00000000;
             1545:out <= 32'h00000000;
             1546:out <= 32'h00000000;
             1547:out <= 32'h00000000;
             1548:out <= 32'h00000000;
             1549:out <= 32'h00000000;
             1550:out <= 32'h00000000;
             1551:out <= 32'h00000000;
             1552:out <= 32'h00000000;
             1553:out <= 32'h00000000;
             1554:out <= 32'h00000000;
             1555:out <= 32'h00000000;
             1556:out <= 32'h00000000;
             1557:out <= 32'h00000000;
             1558:out <= 32'h00000000;
             1559:out <= 32'h00000000;
             1560:out <= 32'h00000000;
             1561:out <= 32'h00000000;
             1562:out <= 32'h00000000;
             1563:out <= 32'h00000000;
             1564:out <= 32'h00000000;
             1565:out <= 32'h00000000;
             1566:out <= 32'h00000000;
             1567:out <= 32'h00000000;
             1568:out <= 32'h00000000;
             1569:out <= 32'h00000000;
             1570:out <= 32'h00000000;
             1571:out <= 32'h00000000;
             1572:out <= 32'h00000000;
             1573:out <= 32'h00000000;
             1574:out <= 32'h00000000;
             1575:out <= 32'h00000000;
             1576:out <= 32'h00000000;
             1577:out <= 32'h00000000;
             1578:out <= 32'h00000000;
             1579:out <= 32'h00000000;
             1580:out <= 32'h00000000;
             1581:out <= 32'h00000000;
             1582:out <= 32'h00000000;
             1583:out <= 32'h00000000;
             1584:out <= 32'h00000000;
             1585:out <= 32'h00000000;
             1586:out <= 32'h00000000;
             1587:out <= 32'h00000000;
             1588:out <= 32'h00000000;
             1589:out <= 32'h00000000;
             1590:out <= 32'h00000000;
             1591:out <= 32'h00000000;
             1592:out <= 32'h00000000;
             1593:out <= 32'h00000000;
             1594:out <= 32'h00000000;
             1595:out <= 32'h00000000;
             1596:out <= 32'h00000000;
             1597:out <= 32'h00000000;
             1598:out <= 32'h00000000;
             1599:out <= 32'h00000000;
             1600:out <= 32'h00000000;
             1601:out <= 32'h00000000;
             1602:out <= 32'h00000000;
             1603:out <= 32'h00000000;
             1604:out <= 32'h00000000;
             1605:out <= 32'h00000000;
             1606:out <= 32'h00000000;
             1607:out <= 32'h00000000;
             1608:out <= 32'h00000000;
             1609:out <= 32'h00000000;
             1610:out <= 32'h00000000;
             1611:out <= 32'h00000000;
             1612:out <= 32'h00000000;
             1613:out <= 32'h00000000;
             1614:out <= 32'h00000000;
             1615:out <= 32'h00000000;
             1616:out <= 32'h00000000;
             1617:out <= 32'h00000000;
             1618:out <= 32'h00000000;
             1619:out <= 32'h00000000;
             1620:out <= 32'h00000000;
             1621:out <= 32'h00000000;
             1622:out <= 32'h00000000;
             1623:out <= 32'h00000000;
             1624:out <= 32'h00000000;
             1625:out <= 32'h00000000;
             1626:out <= 32'h00000000;
             1627:out <= 32'h00000000;
             1628:out <= 32'h00000000;
             1629:out <= 32'h00000000;
             1630:out <= 32'h00000000;
             1631:out <= 32'h00000000;
             1632:out <= 32'h00000000;
             1633:out <= 32'h00000000;
             1634:out <= 32'h00000000;
             1635:out <= 32'h00000000;
             1636:out <= 32'h00000000;
             1637:out <= 32'h00000000;
             1638:out <= 32'h00000000;
             1639:out <= 32'h00000000;
             1640:out <= 32'h00000000;
             1641:out <= 32'h00000000;
             1642:out <= 32'h00000000;
             1643:out <= 32'h00000000;
             1644:out <= 32'h00000000;
             1645:out <= 32'h00000000;
             1646:out <= 32'h00000000;
             1647:out <= 32'h00000000;
             1648:out <= 32'h00000000;
             1649:out <= 32'h00000000;
             1650:out <= 32'h00000000;
             1651:out <= 32'h00000000;
             1652:out <= 32'h00000000;
             1653:out <= 32'h00000000;
             1654:out <= 32'h00000000;
             1655:out <= 32'h00000000;
             1656:out <= 32'h00000000;
             1657:out <= 32'h00000000;
             1658:out <= 32'h00000000;
             1659:out <= 32'h00000000;
             1660:out <= 32'h00000000;
             1661:out <= 32'h00000000;
             1662:out <= 32'h00000000;
             1663:out <= 32'h00000000;
             1664:out <= 32'h00000000;
             1665:out <= 32'h00000000;
             1666:out <= 32'h00000000;
             1667:out <= 32'h00000000;
             1668:out <= 32'h00000000;
             1669:out <= 32'h00000000;
             1670:out <= 32'h00000000;
             1671:out <= 32'h00000000;
             1672:out <= 32'h00000000;
             1673:out <= 32'h00000000;
             1674:out <= 32'h00000000;
             1675:out <= 32'h00000000;
             1676:out <= 32'h00000000;
             1677:out <= 32'h00000000;
             1678:out <= 32'h00000000;
             1679:out <= 32'h00000000;
             1680:out <= 32'h00000000;
             1681:out <= 32'h00000000;
             1682:out <= 32'h00000000;
             1683:out <= 32'h00000000;
             1684:out <= 32'h00000000;
             1685:out <= 32'h00000000;
             1686:out <= 32'h00000000;
             1687:out <= 32'h00000000;
             1688:out <= 32'h00000000;
             1689:out <= 32'h00000000;
             1690:out <= 32'h00000000;
             1691:out <= 32'h00000000;
             1692:out <= 32'h00000000;
             1693:out <= 32'h00000000;
             1694:out <= 32'h00000000;
             1695:out <= 32'h00000000;
             1696:out <= 32'h00000000;
             1697:out <= 32'h00000000;
             1698:out <= 32'h00000000;
             1699:out <= 32'h00000000;
             1700:out <= 32'h00000000;
             1701:out <= 32'h00000000;
             1702:out <= 32'h00000000;
             1703:out <= 32'h00000000;
             1704:out <= 32'h00000000;
             1705:out <= 32'h00000000;
             1706:out <= 32'h00000000;
             1707:out <= 32'h00000000;
             1708:out <= 32'h00000000;
             1709:out <= 32'h00000000;
             1710:out <= 32'h00000000;
             1711:out <= 32'h00000000;
             1712:out <= 32'h00000000;
             1713:out <= 32'h00000000;
             1714:out <= 32'h00000000;
             1715:out <= 32'h00000000;
             1716:out <= 32'h00000000;
             1717:out <= 32'h00000000;
             1718:out <= 32'h00000000;
             1719:out <= 32'h00000000;
             1720:out <= 32'h00000000;
             1721:out <= 32'h00000000;
             1722:out <= 32'h00000000;
             1723:out <= 32'h00000000;
             1724:out <= 32'h00000000;
             1725:out <= 32'h00000000;
             1726:out <= 32'h00000000;
             1727:out <= 32'h00000000;
             1728:out <= 32'h00000000;
             1729:out <= 32'h00000000;
             1730:out <= 32'h00000000;
             1731:out <= 32'h00000000;
             1732:out <= 32'h00000000;
             1733:out <= 32'h00000000;
             1734:out <= 32'h00000000;
             1735:out <= 32'h00000000;
             1736:out <= 32'h00000000;
             1737:out <= 32'h00000000;
             1738:out <= 32'h00000000;
             1739:out <= 32'h00000000;
             1740:out <= 32'h00000000;
             1741:out <= 32'h00000000;
             1742:out <= 32'h00000000;
             1743:out <= 32'h00000000;
             1744:out <= 32'h00000000;
             1745:out <= 32'h00000000;
             1746:out <= 32'h00000000;
             1747:out <= 32'h00000000;
             1748:out <= 32'h00000000;
             1749:out <= 32'h00000000;
             1750:out <= 32'h00000000;
             1751:out <= 32'h00000000;
             1752:out <= 32'h00000000;
             1753:out <= 32'h00000000;
             1754:out <= 32'h00000000;
             1755:out <= 32'h00000000;
             1756:out <= 32'h00000000;
             1757:out <= 32'h00000000;
             1758:out <= 32'h00000000;
             1759:out <= 32'h00000000;
             1760:out <= 32'h00000000;
             1761:out <= 32'h00000000;
             1762:out <= 32'h00000000;
             1763:out <= 32'h00000000;
             1764:out <= 32'h00000000;
             1765:out <= 32'h00000000;
             1766:out <= 32'h00000000;
             1767:out <= 32'h00000000;
             1768:out <= 32'h00000000;
             1769:out <= 32'h00000000;
             1770:out <= 32'h00000000;
             1771:out <= 32'h00000000;
             1772:out <= 32'h00000000;
             1773:out <= 32'h00000000;
             1774:out <= 32'h00000000;
             1775:out <= 32'h00000000;
             1776:out <= 32'h00000000;
             1777:out <= 32'h00000000;
             1778:out <= 32'h00000000;
             1779:out <= 32'h00000000;
             1780:out <= 32'h00000000;
             1781:out <= 32'h00000000;
             1782:out <= 32'h00000000;
             1783:out <= 32'h00000000;
             1784:out <= 32'h00000000;
             1785:out <= 32'h00000000;
             1786:out <= 32'h00000000;
             1787:out <= 32'h00000000;
             1788:out <= 32'h00000000;
             1789:out <= 32'h00000000;
             1790:out <= 32'h00000000;
             1791:out <= 32'h00000000;
             1792:out <= 32'h00000000;
             1793:out <= 32'h00000000;
             1794:out <= 32'h00000000;
             1795:out <= 32'h00000000;
             1796:out <= 32'h00000000;
             1797:out <= 32'h00000000;
             1798:out <= 32'h00000000;
             1799:out <= 32'h00000000;
             1800:out <= 32'h00000000;
             1801:out <= 32'h00000000;
             1802:out <= 32'h00000000;
             1803:out <= 32'h00000000;
             1804:out <= 32'h00000000;
             1805:out <= 32'h00000000;
             1806:out <= 32'h00000000;
             1807:out <= 32'h00000000;
             1808:out <= 32'h00000000;
             1809:out <= 32'h00000000;
             1810:out <= 32'h00000000;
             1811:out <= 32'h00000000;
             1812:out <= 32'h00000000;
             1813:out <= 32'h00000000;
             1814:out <= 32'h00000000;
             1815:out <= 32'h00000000;
             1816:out <= 32'h00000000;
             1817:out <= 32'h00000000;
             1818:out <= 32'h00000000;
             1819:out <= 32'h00000000;
             1820:out <= 32'h00000000;
             1821:out <= 32'h00000000;
             1822:out <= 32'h00000000;
             1823:out <= 32'h00000000;
             1824:out <= 32'h00000000;
             1825:out <= 32'h00000000;
             1826:out <= 32'h00000000;
             1827:out <= 32'h00000000;
             1828:out <= 32'h00000000;
             1829:out <= 32'h00000000;
             1830:out <= 32'h00000000;
             1831:out <= 32'h00000000;
             1832:out <= 32'h00000000;
             1833:out <= 32'h00000000;
             1834:out <= 32'h00000000;
             1835:out <= 32'h00000000;
             1836:out <= 32'h00000000;
             1837:out <= 32'h00000000;
             1838:out <= 32'h00000000;
             1839:out <= 32'h00000000;
             1840:out <= 32'h00000000;
             1841:out <= 32'h00000000;
             1842:out <= 32'h00000000;
             1843:out <= 32'h00000000;
             1844:out <= 32'h00000000;
             1845:out <= 32'h00000000;
             1846:out <= 32'h00000000;
             1847:out <= 32'h00000000;
             1848:out <= 32'h00000000;
             1849:out <= 32'h00000000;
             1850:out <= 32'h00000000;
             1851:out <= 32'h00000000;
             1852:out <= 32'h00000000;
             1853:out <= 32'h00000000;
             1854:out <= 32'h00000000;
             1855:out <= 32'h00000000;
             1856:out <= 32'h00000000;
             1857:out <= 32'h00000000;
             1858:out <= 32'h00000000;
             1859:out <= 32'h00000000;
             1860:out <= 32'h00000000;
             1861:out <= 32'h00000000;
             1862:out <= 32'h00000000;
             1863:out <= 32'h00000000;
             1864:out <= 32'h00000000;
             1865:out <= 32'h00000000;
             1866:out <= 32'h00000000;
             1867:out <= 32'h00000000;
             1868:out <= 32'h00000000;
             1869:out <= 32'h00000000;
             1870:out <= 32'h00000000;
             1871:out <= 32'h00000000;
             1872:out <= 32'h00000000;
             1873:out <= 32'h00000000;
             1874:out <= 32'h00000000;
             1875:out <= 32'h00000000;
             1876:out <= 32'h00000000;
             1877:out <= 32'h00000000;
             1878:out <= 32'h00000000;
             1879:out <= 32'h00000000;
             1880:out <= 32'h00000000;
             1881:out <= 32'h00000000;
             1882:out <= 32'h00000000;
             1883:out <= 32'h00000000;
             1884:out <= 32'h00000000;
             1885:out <= 32'h00000000;
             1886:out <= 32'h00000000;
             1887:out <= 32'h00000000;
             1888:out <= 32'h00000000;
             1889:out <= 32'h00000000;
             1890:out <= 32'h00000000;
             1891:out <= 32'h00000000;
             1892:out <= 32'h00000000;
             1893:out <= 32'h00000000;
             1894:out <= 32'h00000000;
             1895:out <= 32'h00000000;
             1896:out <= 32'h00000000;
             1897:out <= 32'h00000000;
             1898:out <= 32'h00000000;
             1899:out <= 32'h00000000;
             1900:out <= 32'h00000000;
             1901:out <= 32'h00000000;
             1902:out <= 32'h00000000;
             1903:out <= 32'h00000000;
             1904:out <= 32'h00000000;
             1905:out <= 32'h00000000;
             1906:out <= 32'h00000000;
             1907:out <= 32'h00000000;
             1908:out <= 32'h00000000;
             1909:out <= 32'h00000000;
             1910:out <= 32'h00000000;
             1911:out <= 32'h00000000;
             1912:out <= 32'h00000000;
             1913:out <= 32'h00000000;
             1914:out <= 32'h00000000;
             1915:out <= 32'h00000000;
             1916:out <= 32'h00000000;
             1917:out <= 32'h00000000;
             1918:out <= 32'h00000000;
             1919:out <= 32'h00000000;
             1920:out <= 32'h00000000;
             1921:out <= 32'h00000000;
             1922:out <= 32'h00000000;
             1923:out <= 32'h00000000;
             1924:out <= 32'h00000000;
             1925:out <= 32'h00000000;
             1926:out <= 32'h00000000;
             1927:out <= 32'h00000000;
             1928:out <= 32'h00000000;
             1929:out <= 32'h00000000;
             1930:out <= 32'h00000000;
             1931:out <= 32'h00000000;
             1932:out <= 32'h00000000;
             1933:out <= 32'h00000000;
             1934:out <= 32'h00000000;
             1935:out <= 32'h00000000;
             1936:out <= 32'h00000000;
             1937:out <= 32'h00000000;
             1938:out <= 32'h00000000;
             1939:out <= 32'h00000000;
             1940:out <= 32'h00000000;
             1941:out <= 32'h00000000;
             1942:out <= 32'h00000000;
             1943:out <= 32'h00000000;
             1944:out <= 32'h00000000;
             1945:out <= 32'h00000000;
             1946:out <= 32'h00000000;
             1947:out <= 32'h00000000;
             1948:out <= 32'h00000000;
             1949:out <= 32'h00000000;
             1950:out <= 32'h00000000;
             1951:out <= 32'h00000000;
             1952:out <= 32'h00000000;
             1953:out <= 32'h00000000;
             1954:out <= 32'h00000000;
             1955:out <= 32'h00000000;
             1956:out <= 32'h00000000;
             1957:out <= 32'h00000000;
             1958:out <= 32'h00000000;
             1959:out <= 32'h00000000;
             1960:out <= 32'h00000000;
             1961:out <= 32'h00000000;
             1962:out <= 32'h00000000;
             1963:out <= 32'h00000000;
             1964:out <= 32'h00000000;
             1965:out <= 32'h00000000;
             1966:out <= 32'h00000000;
             1967:out <= 32'h00000000;
             1968:out <= 32'h00000000;
             1969:out <= 32'h00000000;
             1970:out <= 32'h00000000;
             1971:out <= 32'h00000000;
             1972:out <= 32'h00000000;
             1973:out <= 32'h00000000;
             1974:out <= 32'h00000000;
             1975:out <= 32'h00000000;
             1976:out <= 32'h00000000;
             1977:out <= 32'h00000000;
             1978:out <= 32'h00000000;
             1979:out <= 32'h00000000;
             1980:out <= 32'h00000000;
             1981:out <= 32'h00000000;
             1982:out <= 32'h00000000;
             1983:out <= 32'h00000000;
             1984:out <= 32'h00000000;
             1985:out <= 32'h00000000;
             1986:out <= 32'h00000000;
             1987:out <= 32'h00000000;
             1988:out <= 32'h00000000;
             1989:out <= 32'h00000000;
             1990:out <= 32'h00000000;
             1991:out <= 32'h00000000;
             1992:out <= 32'h00000000;
             1993:out <= 32'h00000000;
             1994:out <= 32'h00000000;
             1995:out <= 32'h00000000;
             1996:out <= 32'h00000000;
             1997:out <= 32'h00000000;
             1998:out <= 32'h00000000;
             1999:out <= 32'h00000000;
             2000:out <= 32'h00000000;
             2001:out <= 32'h00000000;
             2002:out <= 32'h00000000;
             2003:out <= 32'h00000000;
             2004:out <= 32'h00000000;
             2005:out <= 32'h00000000;
             2006:out <= 32'h00000000;
             2007:out <= 32'h00000000;
             2008:out <= 32'h00000000;
             2009:out <= 32'h00000000;
             2010:out <= 32'h00000000;
             2011:out <= 32'h00000000;
             2012:out <= 32'h00000000;
             2013:out <= 32'h00000000;
             2014:out <= 32'h00000000;
             2015:out <= 32'h00000000;
             2016:out <= 32'h00000000;
             2017:out <= 32'h00000000;
             2018:out <= 32'h00000000;
             2019:out <= 32'h00000000;
             2020:out <= 32'h00000000;
             2021:out <= 32'h00000000;
             2022:out <= 32'h00000000;
             2023:out <= 32'h00000000;
             2024:out <= 32'h00000000;
             2025:out <= 32'h00000000;
             2026:out <= 32'h00000000;
             2027:out <= 32'h00000000;
             2028:out <= 32'h00000000;
             2029:out <= 32'h00000000;
             2030:out <= 32'h00000000;
             2031:out <= 32'h00000000;
             2032:out <= 32'h00000000;
             2033:out <= 32'h00000000;
             2034:out <= 32'h00000000;
             2035:out <= 32'h00000000;
             2036:out <= 32'h00000000;
             2037:out <= 32'h00000000;
             2038:out <= 32'h00000000;
             2039:out <= 32'h00000000;
             2040:out <= 32'h00000000;
             2041:out <= 32'h00000000;
             2042:out <= 32'h00000000;
             2043:out <= 32'h00000000;
             2044:out <= 32'h00000000;
             2045:out <= 32'h00000000;
             2046:out <= 32'h00000000;
             2047:out <= 32'h00000000;

	  endcase
    end
  end

  assign q = oe ? out : 32'bZ;

endmodule

