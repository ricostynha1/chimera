// This program was cloned from: https://github.com/bunny965/yolov5-fpga-hardware-acceleration
// License: GNU General Public License v3.0

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/05/04 00:36:49
// Design Name: 
// Module Name: CSP2_1_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module CSP2_1_tb();
parameter DATA_WIDTH = 16;
parameter D = 3; //Depth of image and filter
parameter H = 4; //Height of image
parameter W = 4; //Width of image
parameter F = 3; //Size of filter
//cbs11
parameter cbs11_K = 2; //Number of filters applied
localparam cbs11_size = cbs11_K*(H-F+1)*(W-F+1);
parameter cbs11_beta =16'b0000000000000000;//0
parameter cbs11_gama = 16'b0011110000000000;//1
parameter cbs11_quarter = 16'b0011010000000000;//1/size
parameter cbs11_channel = cbs11_K;
localparam cbs11_size_div_channel = cbs11_size/cbs11_channel;
//cbs2
parameter cbs2_K = 2; //Number of filters applied
localparam cbs2_size = cbs2_K*(H-F+1)*(W-F+1);
parameter cbs2_beta =16'b0000000000000000;//0
parameter cbs2_gama = 16'b0011110000000000;//1
parameter cbs2_quarter = 16'b0011010000000000;//1/size
localparam cbs2_channel = cbs2_K;
localparam cbs2_size_div_channel = cbs2_size/cbs2_channel;

//cbs12 and cbs13
localparam cbs12_D = cbs11_K; //Depth of image and filter
localparam cbs12_H = (H-F+1); //Height of image
localparam cbs12_W = (W-F+1); //Width of image
localparam cbs12_F = 1; //Number of filters applied
parameter cbs12_K = 2; //Number of filters applied
localparam cbs12_size = cbs12_K*(cbs12_H-cbs12_F+1)*(cbs12_W-cbs12_F+1);
parameter cbs12_beta =16'b0000000000000000;//0
parameter cbs12_gama = 16'b0011110000000000;//1
parameter cbs12_quarter = 16'b0011010000000000;//1/size
localparam cbs12_channel = cbs12_K;
localparam cbs12_size_div_channel = cbs12_size/cbs12_channel;

localparam cbs13_D = cbs12_K; //Depth of image and filter
localparam cbs13_H = (cbs12_H-cbs12_F+3); //Height of image
localparam cbs13_W = (cbs12_W-cbs12_F+3); //Width of image
localparam cbs13_F = 3; //Number of filters applied
parameter cbs13_K = 3; //Number of filters applied
localparam cbs13_size = cbs13_K*(cbs13_H-cbs13_F+1)*(cbs13_W-cbs13_F+1);
parameter cbs13_beta =16'b0000000000000000;//0
parameter cbs13_gama = 16'b0011110000000000;//1
parameter cbs13_quarter = 16'b0011010000000000;//1/size
localparam cbs13_channel = cbs13_K;
localparam cbs13_size_div_channel = cbs13_size/cbs13_channel;


localparam cbso_D = (cbs13_K+cbs2_K); //Depth of image and filter
localparam cbso_H = (H-F+1); //Height of image
localparam cbso_W = (W-F+1); //Width of image
parameter cbso_F = 1; //Size of filter
parameter cbso_K = 2; //Number of filters applied
localparam cbso_size = cbso_K*(cbso_H-cbso_F+1)*(cbso_W-cbso_F+1);
parameter cbso_beta =16'b0000000000000000;//0
parameter cbso_gama = 16'b0011110000000000;//1
parameter cbso_quarter = 16'b0011010000000000;//1/size
localparam cbso_channel = cbso_K;
localparam cbso_size_div_channel = cbso_size/cbso_channel;

reg clk, reset;
reg [D*H*W*DATA_WIDTH-1:0] x;
reg [cbs11_K*D*F*F*DATA_WIDTH-1:0] cbs11_filters;
reg [cbs2_K*D*F*F*DATA_WIDTH-1:0] cbs2_filters;
reg [cbso_K*cbso_D*cbso_F*cbso_F*DATA_WIDTH-1:0] cbso_filters;
reg [cbs12_K*cbs12_D*cbs12_F*cbs12_F*DATA_WIDTH-1:0] cbs12_filters;
reg [cbs13_K*cbs13_D*cbs13_F*cbs13_F*DATA_WIDTH-1:0] cbs13_filters;
wire [DATA_WIDTH*cbso_size-1:0] out;
localparam PERIOD = 100;
integer i;
always #(PERIOD/2) clk = ~clk;
initial begin
#0 reset <=1'b1;
clk<=1'b0;
cbs11_filters<=864'b001111110101110111101010100010100111010011000000011101011101110111110010010101100111000110100111011000010010011011110110010000110000000101100110100110100001100100010000001111100011100101011011011100010101101110101010001000001001011000100011011100010000101000000101010001100110011000000000001001110011100111010111110110110111101010001110100100111110010010001110001111100101111010100111101000110010100101010111111000111101110100111110111010011110011001110111011110010010001111001010100101101011000100000101111011010010100001001100110001001010001101110101001011010110100111010000111100001100011011011011111101011110111101111111111111100101101100001100011110011000100000001110000001000101111010011111000000110100101101001100010110100011010011001100111110111111101111101110111111001010100110101100100111101000001010101111011111001100010100010010100000110111100100101101;
    cbs2_filters<=864'b101111111111111110010101001101000101011100000101111101110001011000001000011011111100010011100100110101001111001111011111111000000110111010111011101001001101001100111001100000111010101001110000010001000111100111100010110101001001000110100011011110010111110110010101000111010000110111111100101101011011111110110000011110100110100010111111001011000010111111001100000110001100010001111101001011010001011011111101001110100110101011110111001101110001110010010001111110000111001011011111000100111110110101000000001110110101010001111100110101101000011001111101011000010001001011010011110111100001101000101000101101011110111010000010011011101101010101001100101000101001101100010011000000111100010100010101000001110001101001101001000001000110100000010110111011000101111110110011100001010011100011111110011110011100010011100001101001000011000000001110000110011010111111111111;
    cbso_filters<=160'b1100100110111101101111001100110100110000100110011010001100011110000111101000111001011111111001001101010111001110101111110001110010011011011111100011111111010010;
    cbs12_filters<=64'b1011111100100010100001011100001000110101110001100101000101011000;
    cbs13_filters<=576'b000011101000000100000100001011010101000100001001001000001000100000100001100011110111000100011011110111101001101001101110111000111010001100011001001110101000010010010110111000111001111100111000001100000010110001110000100000010001001100010101010011100011001011100001110101000000011101001110110001101111111001101100100111101111101010001011011010110101101001100110111011000100100110101100100101011110001011111110111001100000100000110110011110011111100101000001001110011000111010110011101010100100011101111011110100000010111111000100101101111100010011110011110011010110011011011001;
    x<=768'b100000001000111000010100000011100001001010100110101110100100111011000001010000001100110001110010000000010010001011011100011100101110101111100100101111101000000110101000001101010011101000000000101101000111011111111110011000000010010100101110110000110000010001011111000011101110001001111101010010101110110110101101001100100011100011101110001100011001000000111101111010000000001110001010001010001100001110110010111100111000001110111011110000001011100000010101110001010100010011101011000011011011111000111011110010101000101010111001111111100100101011001110110000011100011100001100011101110101011100010001011000111110101001001011001001011011100010000100000011101101011101101000000111000110001000001101100000101101101110001110110110101110110100000100101110110000010100111011;
   # (PERIOD/2) reset<=1'b0;
   #(100*PERIOD)
    for(i=0;i<cbso_size;i=i+1) $display("%b ",out[i*DATA_WIDTH +: DATA_WIDTH]);
    $finish;
end
CSP2_1 UUT (clk,reset,x,cbs11_filters,cbs12_filters,cbs13_filters,cbs2_filters,cbso_filters,out);
endmodule
