// This program was cloned from: https://github.com/lnis-uofu/OpenFPGA
// License: MIT License

module decoder128(datain,dataout);

input [6:0] datain;
output [127:0] dataout;
reg [127:0] dataout;

always @(datain)

begin

	case (datain)
	
		7'b0000000: dataout  <=  128'h00000000000000000000000000000001;
		7'b0000001: dataout  <=  128'h00000000000000000000000000000002;
		7'b0000010: dataout  <=  128'h00000000000000000000000000000004;
		7'b0000011: dataout  <=  128'h00000000000000000000000000000008;
		7'b0000100: dataout  <=  128'h00000000000000000000000000000010;
		7'b0000101: dataout  <=  128'h00000000000000000000000000000020;
		7'b0000110: dataout  <=  128'h00000000000000000000000000000040;
		7'b0000111: dataout	 <=  128'h00000000000000000000000000000080;
		7'b0001000: dataout  <=  128'h00000000000000000000000000000100;
		7'b0001001: dataout  <=  128'h00000000000000000000000000000200;
		7'b0001010: dataout  <=  128'h00000000000000000000000000000400;
		7'b0001011: dataout  <=  128'h00000000000000000000000000000800;
		7'b0001100: dataout  <=  128'h00000000000000000000000000001000;
		7'b0001101: dataout  <=  128'h00000000000000000000000000002000;
		7'b0001110: dataout  <=  128'h00000000000000000000000000004000;
		7'b0001111: dataout	 <=  128'h00000000000000000000000000008000; 		
    7'b0010000: dataout  <=  128'h00000000000000000000000000010000;
		7'b0010001: dataout  <=  128'h00000000000000000000000000020000;
		7'b0010010: dataout  <=  128'h00000000000000000000000000040000;
		7'b0010011: dataout  <=  128'h00000000000000000000000000080000;
		7'b0010100: dataout  <=  128'h00000000000000000000000000100000;
		7'b0010101: dataout  <=  128'h00000000000000000000000000200000;
		7'b0010110: dataout  <=  128'h00000000000000000000000000400000;
		7'b0010111: dataout  <=  128'h00000000000000000000000000800000;
		7'b0011000: dataout	 <=  128'h00000000000000000000000001000000;
		7'b0011001: dataout  <=  128'h00000000000000000000000002000000;
		7'b0011010: dataout  <=  128'h00000000000000000000000004000000;
		7'b0011011: dataout  <=  128'h00000000000000000000000008000000;
		7'b0011100: dataout  <=  128'h00000000000000000000000010000000;
		7'b0011101: dataout  <=  128'h00000000000000000000000020000000;
		7'b0011110: dataout  <=  128'h00000000000000000000000040000000;
		7'b0011111: dataout  <=  128'h00000000000000000000000080000000;                                        
	  7'b0100000: dataout  <=  128'h00000000000000000000000100000000;                  
	  7'b0100001: dataout  <=  128'h00000000000000000000000200000000;
	  7'b0100010: dataout  <=  128'h00000000000000000000000400000000;
	  7'b0100011: dataout  <=  128'h00000000000000000000000800000000;
	  7'b0100100: dataout  <=  128'h00000000000000000000001000000000;
	  7'b0100101: dataout  <=  128'h00000000000000000000002000000000;
	  7'b0100110: dataout  <=  128'h00000000000000000000004000000000;
	  7'b0100111: dataout  <=  128'h00000000000000000000008000000000;
	  7'b0101000: dataout  <=  128'h00000000000000000000010000000000;
	  7'b0101001: dataout  <=  128'h00000000000000000000020000000000;
	  7'b0101010: dataout  <=  128'h00000000000000000000040000000000;
	  7'b0101011: dataout  <=  128'h00000000000000000000080000000000;
	  7'b0101100: dataout  <=  128'h00000000000000000000100000000000;
	  7'b0101101: dataout  <=  128'h00000000000000000000200000000000;
	  7'b0101110: dataout  <=  128'h00000000000000000000400000000000;
	  7'b0101111: dataout  <=  128'h00000000000000000000800000000000;                                                                  
	  7'b0110000: dataout  <=  128'h00000000000000000001000000000000;
	  7'b0110001: dataout  <=  128'h00000000000000000002000000000000;
	  7'b0110010: dataout  <=  128'h00000000000000000004000000000000;
	  7'b0110011: dataout  <=  128'h00000000000000000008000000000000;
	  7'b0110100: dataout  <=  128'h00000000000000000010000000000000;
	  7'b0110101: dataout  <=  128'h00000000000000000020000000000000;
	  7'b0110110: dataout  <=  128'h00000000000000000040000000000000;
	  7'b0110111: dataout  <=  128'h00000000000000000080000000000000;
	  7'b0111000: dataout  <=  128'h00000000000000000100000000000000;
	  7'b0111001: dataout  <=  128'h00000000000000000200000000000000;
	  7'b0111010: dataout  <=  128'h00000000000000000400000000000000;
	  7'b0111011: dataout  <=  128'h00000000000000000800000000000000;
	  7'b0111100: dataout  <=  128'h00000000000000001000000000000000;                  
	  7'b0111101: dataout  <=  128'h00000000000000002000000000000000;                  
	  7'b0111110: dataout  <=  128'h00000000000000004000000000000000;                  
	  7'b0111111: dataout  <=  128'h00000000000000008000000000000000;                  
	  7'b1000000: dataout  <=  128'h00000000000000010000000000000000;                   
	  7'b1000001: dataout  <=  128'h00000000000000020000000000000000;                   
	  7'b1000010: dataout  <=  128'h00000000000000040000000000000000;
    7'b1000011: dataout  <=  128'h00000000000000080000000000000000;
    7'b1000100: dataout  <=  128'h00000000000000100000000000000000;
    7'b1000101: dataout  <=  128'h00000000000000200000000000000000;
    7'b1000110: dataout  <=  128'h00000000000000400000000000000000;
    7'b1000111: dataout  <=  128'h00000000000000800000000000000000;
    7'b1001000: dataout  <=  128'h00000000000001000000000000000000;
    7'b1001001: dataout  <=  128'h00000000000002000000000000000000;
    7'b1001010: dataout  <=  128'h00000000000004000000000000000000;
    7'b1001011: dataout  <=  128'h00000000000008000000000000000000;
    7'b1001100: dataout  <=  128'h00000000000010000000000000000000;
    7'b1001101: dataout  <=  128'h00000000000020000000000000000000;
    7'b1001110: dataout  <=  128'h00000000000040000000000000000000;
    7'b1001111: dataout  <=  128'h00000000000080000000000000000000;
    7'b1010000: dataout  <=  128'h00000000000100000000000000000000;
    7'b1010001: dataout  <=  128'h00000000000200000000000000000000;
    7'b1010010: dataout  <=  128'h00000000000400000000000000000000;
    7'b1010011: dataout  <=  128'h00000000000800000000000000000000;
    7'b1010100: dataout  <=  128'h00000000001000000000000000000000;
    7'b1010101: dataout  <=  128'h00000000002000000000000000000000;
    7'b1010110: dataout  <=  128'h00000000004000000000000000000000;
    7'b1010111: dataout  <=  128'h00000000008000000000000000000000;
    7'b1011000: dataout  <=  128'h00000000010000000000000000000000;
    7'b1011001: dataout  <=  128'h00000000020000000000000000000000;
    7'b1011010: dataout  <=  128'h00000000040000000000000000000000;
    7'b1011011: dataout  <=  128'h00000000080000000000000000000000;
    7'b1011100: dataout  <=  128'h00000000100000000000000000000000;
    7'b1011101: dataout  <=  128'h00000000200000000000000000000000;
    7'b1011110: dataout  <=  128'h00000000400000000000000000000000;
    7'b1011111: dataout  <=  128'h00000000800000000000000000000000;
    7'b1100000: dataout  <=  128'h00000001000000000000000000000000;
    7'b1100001: dataout  <=  128'h00000002000000000000000000000000;
    7'b1100010: dataout  <=  128'h00000004000000000000000000000000;
    7'b1100011: dataout  <=  128'h00000008000000000000000000000000;
    7'b1100100: dataout  <=  128'h00000010000000000000000000000000;
    7'b1100101: dataout  <=  128'h00000020000000000000000000000000;
    7'b1100110: dataout  <=  128'h00000040000000000000000000000000;
    7'b1100111: dataout  <=  128'h00000080000000000000000000000000;
    7'b1101000: dataout  <=  128'h00000100000000000000000000000000;
    7'b1101001: dataout  <=  128'h00000200000000000000000000000000;
    7'b1101010: dataout  <=  128'h00000400000000000000000000000000;
    7'b1101011: dataout  <=  128'h00000800000000000000000000000000;
    7'b1101100: dataout  <=  128'h00001000000000000000000000000000;
    7'b1101101: dataout  <=  128'h00002000000000000000000000000000;
    7'b1101110: dataout  <=  128'h00004000000000000000000000000000;
    7'b1101111: dataout  <=  128'h00008000000000000000000000000000;
    7'b1110000: dataout  <=  128'h00010000000000000000000000000000;
    7'b1110001: dataout  <=  128'h00020000000000000000000000000000;
    7'b1110010: dataout  <=  128'h00040000000000000000000000000000;
    7'b1110011: dataout  <=  128'h00080000000000000000000000000000;
    7'b1110100: dataout  <=  128'h00100000000000000000000000000000;
    7'b1110101: dataout  <=  128'h00200000000000000000000000000000;
    7'b1110110: dataout  <=  128'h00400000000000000000000000000000;
    7'b1110111: dataout  <=  128'h00800000000000000000000000000000;
    7'b1111000: dataout  <=  128'h01000000000000000000000000000000;
    7'b1111001: dataout  <=  128'h02000000000000000000000000000000;
    7'b1111010: dataout  <=  128'h04000000000000000000000000000000;
    7'b1111011: dataout  <=  128'h08000000000000000000000000000000;
    7'b1111100: dataout  <=  128'h10000000000000000000000000000000;
    7'b1111101: dataout  <=  128'h20000000000000000000000000000000;
    7'b1111110: dataout  <=  128'h40000000000000000000000000000000;
    7'b1111111:  dataout  <=  128'h80000000000000000000000000000000;
    
    
    
    default: dataout<=128'h0;
		endcase
end
endmodule
