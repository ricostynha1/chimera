// This program was cloned from: https://github.com/Nilesh002/Multiplication-and-Accumulation-Unit-MAC-
// License: MIT License

module add6(a,b,s);
input [5:0]a,b;
output [5:0]s;

assign s=a+b;


endmodule
