// This program was cloned from: https://github.com/emu-russia/SEGAChips
// License: Creative Commons Zero v1.0 Universal

module ym6045
	(
	input MCLK,
	input MCLK_e,
	input VCLK,
	input ZCLK,
	input VD8_i,
	input [15:7] ZA_i,
	input ZA0_i,
	input [22:7] VA_i,
	input ZRD_i,
	input M1,
	input ZWR_i,
	input BGACK_i,
	input BG,
	input IORQ,
	input RW_i,
	input UDS_i,
	input AS_i,
	input DTACK_i,
	input LDS_i,
	input CAS0,
	input M3,
	input WRES,
	input CART,
	input OE0,
	input WAIT_i,
	input ZBAK,
	input MREQ_i,
	input FC0,
	input FC1,
	input SRES,
	input test_mode_0,
	input ZD0_i,
	input HSYNC,
	output VD8_o,
	output ZA0_o,
	output [15:8] ZA_o,
	output [22:7] VA_o,
	output ZRD_o,
	output UDS_o,
	output ZWR_o,
	output BGACK_o,
	output AS_o,
	output RW_d,
	output RW_o,
	output LDS_o,
	output strobe_dir,
	output DTACK_o,
	output BR,
	output IA14,
	output TIME,
	output CE0,
	output FDWR,
	output FDC,
	output ROM,
	output ASEL,
	output EOE,
	output NOE,
	output RAS2,
	output CAS2,
	output REF,
	output ZRAM,
	output WAIT_o,
	output ZBR,
	output NMI,
	output ZRES,
	output SOUND,
	output VZ,
	output MREQ_o,
	output VRES,
	output VPA,
	output VDPM,
	output IO,
	output ZV,
	output INTAK,
	output EDCLK,
	output vtoz,
	output w12,
	output w131,
	output w142,
	output w310,
	output w353
	);
	
	wire pal_trap = ~1'h1;
	
	wire EDCLK2;
	
	reg edclk_buf;
	
	always @(posedge MCLK)
	begin
		edclk_buf <= EDCLK2;
	end
	
	assign EDCLK = edclk_buf;
	
	assign vtoz = VZ;
	
	ym6045c arb
		(
		.VA8_d(w131),
		.VA21_d(w142),
		.TPAL(~pal_trap),
		.n_LDS_d(strobe_dir),
		
		.VA8_o(VA_o[7]),
		.VA8_i(VA_i[7]),
		.VA9_o(VA_o[8]),
		.VA9_i(VA_i[8]),
		.VA10_o(VA_o[9]),
		.VA10_i(VA_i[9]),
		.VA11_o(VA_o[10]),
		.VA11_i(VA_i[10]),
		.VA12_o(VA_o[11]),
		.VA12_i(VA_i[11]),
		.VA13_o(VA_o[12]),
		.VA13_i(VA_i[12]),
		.VA14_o(VA_o[13]),
		.VA14_i(VA_i[13]),
		.VA15_o(VA_o[14]),
		.VA15_i(VA_i[14]),
		.VA16_o(VA_o[15]),
		.VA16_i(VA_i[15]),
		.VA17_o(VA_o[16]),
		.VA17_i(VA_i[16]),
		.VA18_o(VA_o[17]),
		.VA18_i(VA_i[17]),
		.VA19_o(VA_o[18]),
		.VA19_i(VA_i[18]),
		.VA20_o(VA_o[19]),
		.VA20_i(VA_i[19]),
		.VA21_o(VA_o[20]),
		.VA21_i(VA_i[20]),
		.VA22_o(VA_o[21]),
		.VA22_i(VA_i[21]),
		.VA23_o(VA_o[22]),
		.VA23_i(VA_i[22]),
		.FC0(FC0),
		.FC1(FC1),
		.n_VPA(VPA),
		.n_RESET(VRES),
		.D8_o(VD8_o),
		.D8_d(w12),
		.D8_i(VD8_i),
		.VCLK(VCLK),
		.n_TIME(TIME),
		.n_CAS0(CAS0),
		.n_DTACK_d(DTACK_o),
		.n_DTACK_i(DTACK_i),
		.RW_i(RW_i),
		.RW_d(RW_d),
		.RW_o(RW_o),
		.n_LDS_o(LDS_o),
		.n_LDS_i(LDS_i),
		.n_UDS_o(UDS_o),
		.n_UDS_i(UDS_i),
		.n_AS_o(AS_o),
		.n_AS_i(AS_i),
		.n_INTAK(INTAK),
		.n_VDPM(VDPM),
		.n_BG(BG),
		.n_BGACK_i(BGACK_i),
		.n_BGACK_d(BGACK_o),
		.n_BR(BR),
		.i_EOE(EOE),
		.IA14(IA14),
		.n_NOE(NOE),
		.EDCK(EDCLK2),
		.n_OE0(OE0),
		.n_HSYNC(HSYNC),
		.MCLK(MCLK_e),
		.n_SOUND(SOUND),
		.ZCLK(ZCLK),
		.n_WRES(WRES),
		.n_ZRAM(ZRAM),
		.n_REF(REF),
		.n_M1(M1),
		.n_ZRES(ZRES),
		.n_ZBR(ZBR),
		.n_WAIT_d(WAIT_o),
		.n_WAIT_i(WAIT_i),
		.n_ZBAK(ZBAK),
		.n_ZWR_o(ZWR_o),
		.n_ZWR_i(ZWR_i),
		.n_ZRD_i(ZRD_i),
		.n_ZRD_o(ZRD_o),
		.n_IREQ(IORQ),
		.n_MREQ_i(MREQ_i),
		.n_MREQ_o(MREQ_o),
		.n_NMI(NMI),
		.n_ZA0_i(ZA0_i),
		.n_ZA0_o(ZA0_o),
		.ZA7(ZA_i[7]),
		.ZA8_i(ZA_i[8]),
		.ZA8_o(ZA_o[8]),
		.ZA9_i(ZA_i[9]),
		.ZA9_o(ZA_o[9]),
		.ZA10_i(ZA_i[10]),
		.ZA10_o(ZA_o[10]),
		.ZA11_i(ZA_i[11]),
		.ZA11_o(ZA_o[11]),
		.ZA12_i(ZA_i[12]),
		.ZA12_o(ZA_o[12]),
		.ZA13_i(ZA_i[13]),
		.ZA13_o(ZA_o[13]),
		.ZA14_i(ZA_i[14]),
		.ZA14_o(ZA_o[14]),
		.ZA15_i(ZA_i[15]),
		.ZA15_o(ZA_o[15]),
		.ZD0(ZD0_i),
		.n_FDWR(FDWR),
		.n_FDC(FDC),
		.n_ROM(ROM),
		.n_ASEL(ASEL),
		.n_CAS2(CAS2),
		.n_RAS2(RAS2),
		.n_CE0(CE0),
		.n_VTOZ(VZ),
		.n_ZTOV(ZV),
		.n_SRES(SRES),
		.n_IO(IO),
		.n_M3(M3),
		.n_CART(CART),
		.pin99(w353),
		.pin100(w310)
		);
	
endmodule
