// This program was cloned from: https://github.com/apuder/TRS-IO
// License: GNU General Public License v3.0

//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.9 Beta-4 Education
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Sun Feb 04 09:12:09 2024

module blk_mem_gen_4 (douta, doutb, clka, ocea, cea, reseta, wrea, clkb, oceb, ceb, resetb, wreb, ada, dina, adb, dinb);

output [7:0] douta;
output [7:0] doutb;
input clka;
input ocea;
input cea;
input reseta;
input wrea;
input clkb;
input oceb;
input ceb;
input resetb;
input wreb;
input [14:0] ada;
input [7:0] dina;
input [14:0] adb;
input [7:0] dinb;

wire [14:0] dpb_inst_0_douta_w;
wire [0:0] dpb_inst_0_douta;
wire [14:0] dpb_inst_0_doutb_w;
wire [0:0] dpb_inst_0_doutb;
wire [14:0] dpb_inst_1_douta_w;
wire [1:1] dpb_inst_1_douta;
wire [14:0] dpb_inst_1_doutb_w;
wire [1:1] dpb_inst_1_doutb;
wire [14:0] dpb_inst_2_douta_w;
wire [2:2] dpb_inst_2_douta;
wire [14:0] dpb_inst_2_doutb_w;
wire [2:2] dpb_inst_2_doutb;
wire [14:0] dpb_inst_3_douta_w;
wire [3:3] dpb_inst_3_douta;
wire [14:0] dpb_inst_3_doutb_w;
wire [3:3] dpb_inst_3_doutb;
wire [11:0] dpb_inst_4_douta_w;
wire [3:0] dpb_inst_4_douta;
wire [11:0] dpb_inst_4_doutb_w;
wire [3:0] dpb_inst_4_doutb;
wire [14:0] dpb_inst_5_douta_w;
wire [4:4] dpb_inst_5_douta;
wire [14:0] dpb_inst_5_doutb_w;
wire [4:4] dpb_inst_5_doutb;
wire [14:0] dpb_inst_6_douta_w;
wire [5:5] dpb_inst_6_douta;
wire [14:0] dpb_inst_6_doutb_w;
wire [5:5] dpb_inst_6_doutb;
wire [14:0] dpb_inst_7_douta_w;
wire [6:6] dpb_inst_7_douta;
wire [14:0] dpb_inst_7_doutb_w;
wire [6:6] dpb_inst_7_doutb;
wire [14:0] dpb_inst_8_douta_w;
wire [7:7] dpb_inst_8_douta;
wire [14:0] dpb_inst_8_doutb_w;
wire [7:7] dpb_inst_8_doutb;
wire [11:0] dpb_inst_9_douta_w;
wire [7:4] dpb_inst_9_douta;
wire [11:0] dpb_inst_9_doutb_w;
wire [7:4] dpb_inst_9_doutb;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire cea_w;
wire ceb_w;
wire gw_gnd;

assign cea_w = ~wrea & cea;
assign ceb_w = ~wreb & ceb;
assign gw_gnd = 1'b0;

DPB dpb_inst_0 (
    .DOA({dpb_inst_0_douta_w[14:0],dpb_inst_0_douta[0]}),
    .DOB({dpb_inst_0_doutb_w[14:0],dpb_inst_0_doutb[0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[0]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[0]})
);

defparam dpb_inst_0.READ_MODE0 = 1'b1;
defparam dpb_inst_0.READ_MODE1 = 1'b1;
defparam dpb_inst_0.WRITE_MODE0 = 2'b00;
defparam dpb_inst_0.WRITE_MODE1 = 2'b00;
defparam dpb_inst_0.BIT_WIDTH_0 = 1;
defparam dpb_inst_0.BIT_WIDTH_1 = 1;
defparam dpb_inst_0.BLK_SEL_0 = 3'b000;
defparam dpb_inst_0.BLK_SEL_1 = 3'b000;
defparam dpb_inst_0.RESET_MODE = "SYNC";
defparam dpb_inst_0.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_01 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_03 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_05 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_06 = 256'h0000FFBE303FFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_07 = 256'h0000FFBF203FFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_08 = 256'h0000FFBF303FFFFFFFFF81FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_09 = 256'h0000FFBF383FF0001FFFFFFE1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_0A = 256'h0000FFBF207FE00000000FFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_0B = 256'h0000FFBF307FE08000000001FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_0C = 256'h0000FFBF387FF08000000000FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_0D = 256'h0000FFBF3C7FE08000000000F80000000000000100000000000FFFFFFFFF1FFF;
defparam dpb_inst_0.INIT_RAM_0E = 256'h0000FFBF387FE08001008000FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7F;
defparam dpb_inst_0.INIT_RAM_0F = 256'h0000FFBF3C7FE08001000000FBFFFF000000000000000000000000000000071F;
defparam dpb_inst_0.INIT_RAM_10 = 256'h0000FFBF3C7FE08000000000FBFFF8000000000000000000000000000008001F;
defparam dpb_inst_0.INIT_RAM_11 = 256'h0000FFBF3C7FE08000000C00FBFFF0000000000000000000000000000008001F;
defparam dpb_inst_0.INIT_RAM_12 = 256'h0000FFBF3C7FE08000000000FBFFF0038000000002555555555500000008001F;
defparam dpb_inst_0.INIT_RAM_13 = 256'h0000FFBF3C7FE08000000000FBFFF0007007FFFFFFFFFFFFFFFFFFFF8008004F;
defparam dpb_inst_0.INIT_RAM_14 = 256'h0000FFBF387FE08000140C00FBFFF000087FFFFFFFFFFFFFFFFFFFFFE008004F;
defparam dpb_inst_0.INIT_RAM_15 = 256'h0000FFBF307FE08000000000FBFFF00001FFFFFFFFFFFFFFFFFFFFFFF008004F;
defparam dpb_inst_0.INIT_RAM_16 = 256'h0000FFBF3C7FE08000000000F9FFF00003FFFFFFFFFFFFFFFF03FFFFFC08004F;
defparam dpb_inst_0.INIT_RAM_17 = 256'h0000FFBF387FE08000040000F800700003FFFFFFFFFFFC000023FFFFFC08000F;
defparam dpb_inst_0.INIT_RAM_18 = 256'h0000FFBF347FE08000000000F800300003FFFFFFFFFFFC000023FFFFFC08000F;
defparam dpb_inst_0.INIT_RAM_19 = 256'h0000FFBF3C7FE08000004000F80030000FFFFFFFFFFFFFFFFF03FFFFFE08000F;
defparam dpb_inst_0.INIT_RAM_1A = 256'h0000FFBE387FE08000046000FBFFF0000FFFFFFFFFFFFC000003FFFFFE0C000F;
defparam dpb_inst_0.INIT_RAM_1B = 256'h0000FFBE3C7FE08000000038F80070000FFFFFFFFFFFFC3FFFE3FFFFFE08000F;
defparam dpb_inst_0.INIT_RAM_1C = 256'h0000FFBE3C7FE08000000000F80010001FFFFFFFFFFFFFE01F23FFFFFE04000F;
defparam dpb_inst_0.INIT_RAM_1D = 256'h0000FFBE387FE08000040000F80010001FFFFFFFFFFFFC050043FFFFFE04000F;
defparam dpb_inst_0.INIT_RAM_1E = 256'h0000FFBE3C7FE08001000038F81FF0001FFFFFFFFFFFFC00000FFFFFFE04000F;
defparam dpb_inst_0.INIT_RAM_1F = 256'h0000FFBE3C7FE08000000003F8FFF0001FFFFFFFFFFFFFFFFFFFFFFFFE04002F;
defparam dpb_inst_0.INIT_RAM_20 = 256'h0000FFBE387FE08000040002F80010001FFFFFFFFFFFFC47C003FFFFFE04002F;
defparam dpb_inst_0.INIT_RAM_21 = 256'h0000FFBE3C7FE08001000006F80030001FFFFFFFFFFFF8401021FFFFFF04002F;
defparam dpb_inst_0.INIT_RAM_22 = 256'h0000FFBE3C7FE00000000C0FF80030001FFFFFFFFFFFFC1F0700FFFFFF04002F;
defparam dpb_inst_0.INIT_RAM_23 = 256'h0000FFBE3C7FE00000040002FBFFF8001FFFFFFFFFFFFFE1FFFFFFFFFF04002F;
defparam dpb_inst_0.INIT_RAM_24 = 256'h0000FFBE3C7FE08001000001F80038001FFFFFFFFFFFFFFE27FFFFFFFF07002F;
defparam dpb_inst_0.INIT_RAM_25 = 256'h0000FFBE3C7FE00000000C0FF80018001FFFFFFFFFFFFFFE27FFFFFFFF07002F;
defparam dpb_inst_0.INIT_RAM_26 = 256'h0000FFBE3C7FE00000000003F80038001FFFFFFFFFFFFFFFFFFFFFFFFE07002F;
defparam dpb_inst_0.INIT_RAM_27 = 256'h0000FFBE3C7FE00000000003F807F8041FFFFFFFFFFFFC000003FFFFFE01002F;
defparam dpb_inst_0.INIT_RAM_28 = 256'h0000FFBE3C7FE00000000C0FF87FF8041FFFFFFFFFFFFC000003FFFFFE010C2F;
defparam dpb_inst_0.INIT_RAM_29 = 256'h0000FFBE387FE00000000001F80018041FFFFFFFFFFFFFFE07FFFFFFFE010F2F;
defparam dpb_inst_0.INIT_RAM_2A = 256'h0000FFBE387FE00001000001F80018000FFFFFFFFFFFFF830C0FFFFFFE010FEF;
defparam dpb_inst_0.INIT_RAM_2B = 256'h0000FFBE3C7FE0400000000FF84438040FFFFFFFFFFFFC20F043FFFFFC010FEF;
defparam dpb_inst_0.INIT_RAM_2C = 256'h0000FFBE307FE04000000009FBFFF8000FFFFFFFFFFFF847FF21FFFFFC010FEF;
defparam dpb_inst_0.INIT_RAM_2D = 256'h0000FFBE287FE04001802001F800180003FFFFFFFFFFFC21FC23FFFFFC010FEF;
defparam dpb_inst_0.INIT_RAM_2E = 256'h0000FFBE307FE04000FF4001F800180003FFFFFFFFFFFF860707FFFFFC010FEF;
defparam dpb_inst_0.INIT_RAM_2F = 256'h0000FFBE387FE04000FF001FF800780001FFFFFFFFFFFFFC01FFFFFFF0010FEF;
defparam dpb_inst_0.INIT_RAM_30 = 256'h0000FFBE3C7FE04001FF0000FBFFF80200FFFFFFFFFFFFFFFFFFFFFFE0030FEF;
defparam dpb_inst_0.INIT_RAM_31 = 256'h0000FFBE387FF04001FF0000FBFFF802000FFFFFFFFFFFFFFFFFFFFF80014FEF;
defparam dpb_inst_0.INIT_RAM_32 = 256'h0000FFBE307FE04000FF0010FBFFF80000000000FFFFFFFFFFFC000000014FEF;
defparam dpb_inst_0.INIT_RAM_33 = 256'h0000FFBE307FF04000000800FBFFF80000000000000000000000000000010FEF;
defparam dpb_inst_0.INIT_RAM_34 = 256'h0000FFBE387FF04000040000FBFFF80000000000000000000000000000010FEF;
defparam dpb_inst_0.INIT_RAM_35 = 256'h0000FFBE307FF04000000180FBF3F80000000000000000000000000000010FEF;
defparam dpb_inst_0.INIT_RAM_36 = 256'h0000FFBE207FF04020073800FBC2F80000000000007FFFFFFFFE000000010FEF;
defparam dpb_inst_0.INIT_RAM_37 = 256'h0000FFBE207FF04000000000FBFFF800000000000040003F8183080000010FEF;
defparam dpb_inst_0.INIT_RAM_38 = 256'h0000FFBE207FF04000000000FBFFF800000000000040801D8083000000010BEF;
defparam dpb_inst_0.INIT_RAM_39 = 256'h0000FFBE007FF04000000000FB85F800000000000040881D8081000200010BEF;
defparam dpb_inst_0.INIT_RAM_3A = 256'h0000FFBE287FF0000000C1E0FBC1F800000000000040081F8001000001018FEF;
defparam dpb_inst_0.INIT_RAM_3B = 256'h0000FFBE307FF00004000000FBFFF800000000000040001D8081000000018FEF;
defparam dpb_inst_0.INIT_RAM_3C = 256'h0000FFBE007FF00000000000FBFFF800000000000040001F8081000000018FEF;
defparam dpb_inst_0.INIT_RAM_3D = 256'h0000FFB2007FF0000030C1C0FBFFF80000000000007FFFFFFFFF000000010FFF;
defparam dpb_inst_0.INIT_RAM_3E = 256'h0000FFB2207FF00000000040FBFFF80000000000000000000000000000018FF3;
defparam dpb_inst_0.INIT_RAM_3F = 256'h0000FFBE007FF00020000000FBFFFC0000000000000000000000000000003033;

DPB dpb_inst_1 (
    .DOA({dpb_inst_1_douta_w[14:0],dpb_inst_1_douta[1]}),
    .DOB({dpb_inst_1_doutb_w[14:0],dpb_inst_1_doutb[1]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[1]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[1]})
);

defparam dpb_inst_1.READ_MODE0 = 1'b1;
defparam dpb_inst_1.READ_MODE1 = 1'b1;
defparam dpb_inst_1.WRITE_MODE0 = 2'b00;
defparam dpb_inst_1.WRITE_MODE1 = 2'b00;
defparam dpb_inst_1.BIT_WIDTH_0 = 1;
defparam dpb_inst_1.BIT_WIDTH_1 = 1;
defparam dpb_inst_1.BLK_SEL_0 = 3'b000;
defparam dpb_inst_1.BLK_SEL_1 = 3'b000;
defparam dpb_inst_1.RESET_MODE = "SYNC";
defparam dpb_inst_1.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_01 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_03 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_05 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_06 = 256'h0000FF9E203FF87FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_07 = 256'h0000FFBF303FFFFFE1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_08 = 256'h0000FFBF103FFFFFFFFF87FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_09 = 256'h0000FFBF383FF0001FFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_0A = 256'h0000FFBF207FE00000001FFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_0B = 256'h0000FFBF307FE08000000001FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_0C = 256'h0000FFBF387FE08000000000FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_0D = 256'h0000FFBF3C7FE08000000000FBFFFFFFFFF80000000000000007FFFFFFFF3FFF;
defparam dpb_inst_1.INIT_RAM_0E = 256'h0000FFBF387FE08001008000FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFF;
defparam dpb_inst_1.INIT_RAM_0F = 256'h0000FFBF3C7FE08001000000FBFFFF000000000000000000000000000000071F;
defparam dpb_inst_1.INIT_RAM_10 = 256'h0000FFBF3C7FE08000000018FBFFF8000000000000000000000000000008001F;
defparam dpb_inst_1.INIT_RAM_11 = 256'h0000FFBF3C7FE08000000C00FBFFF0000000000000000000000000000008005F;
defparam dpb_inst_1.INIT_RAM_12 = 256'h0000FFBF387FE08004000000FBFFF0030000000000000000000000000008001F;
defparam dpb_inst_1.INIT_RAM_13 = 256'h0000FFBF3C7FE08000000000FBFFF0007007FFFFFFFFFFFFFFFFFFFF8008004F;
defparam dpb_inst_1.INIT_RAM_14 = 256'h0000FFBF3C7FE08000000C00FBFFF000087FFFFFFFFFFFFFFFFFFFFFE008004F;
defparam dpb_inst_1.INIT_RAM_15 = 256'h0000FFBF387FE08000000000FBFFF00001FFFFFFFFFFFFFFFFFFFFFFF008004F;
defparam dpb_inst_1.INIT_RAM_16 = 256'h0000FFBF387FE08004004000F807F00001FFFFFFFFFFFFFFFF03FFFFF008004F;
defparam dpb_inst_1.INIT_RAM_17 = 256'h0000FFBF387FE08000340000FBFFF00003FFFFFFFFFFFC000023FFFFFC08000F;
defparam dpb_inst_1.INIT_RAM_18 = 256'h0000FFBF307FE08000000000F800700003FFFFFFFFFFFC000023FFFFFC08000F;
defparam dpb_inst_1.INIT_RAM_19 = 256'h0000FFBF3C7FE08000006000F80030000FFFFFFFFFFFFFFFFF03FFFFFE08000F;
defparam dpb_inst_1.INIT_RAM_1A = 256'h0000FFBE3C7FE08000140000F80030000FFFFFFFFFFFFFFFFFFFFFFFFE08000F;
defparam dpb_inst_1.INIT_RAM_1B = 256'h0000FFBE3C7FE08000000010FBFFF0000FFFFFFFFFFFFC7FFFE3FFFFFE08000F;
defparam dpb_inst_1.INIT_RAM_1C = 256'h0000FFBE3C7FE08000000000F80030001FFFFFFFFFFFFFE01F23FFFFFE04000F;
defparam dpb_inst_1.INIT_RAM_1D = 256'h0000FFBE387FE08000040000F80010001FFFFFFFFFFFFC050043FFFFFE04000F;
defparam dpb_inst_1.INIT_RAM_1E = 256'h0000FFBE3C7FE08000000038F80430001FFFFFFFFFFFFC00000FFFFFFE04000F;
defparam dpb_inst_1.INIT_RAM_1F = 256'h0000FFBE3C7FE08000000003F8FFF0001FFFFFFFFFFFFCFFFFFFFFFFFE04000F;
defparam dpb_inst_1.INIT_RAM_20 = 256'h0000FFBE387FE08000040002F801F0001FFFFFFFFFFFFC07E003FFFFFE04002F;
defparam dpb_inst_1.INIT_RAM_21 = 256'h0000FFBE387FE0800100003EF80010001FFFFFFFFFFFF8421021FFFFFF04002F;
defparam dpb_inst_1.INIT_RAM_22 = 256'h0000FFBE3C7FE00000000C07F80030001FFFFFFFFFFFFC0F0701FFFFFF04002F;
defparam dpb_inst_1.INIT_RAM_23 = 256'h0000FFBE3C7FE00000000002F84478001FFFFFFFFFFFFF80FFFFFFFFFF04002F;
defparam dpb_inst_1.INIT_RAM_24 = 256'h0000FFBE3C7FE0000100003EFBFFF8001FFFFFFFFFFFFFFE07FFFFFFFF07002F;
defparam dpb_inst_1.INIT_RAM_25 = 256'h0000FFBE3C7FE0000000000FF80038001FFFFFFFFFFFFFFE27FFFFFFFF07002F;
defparam dpb_inst_1.INIT_RAM_26 = 256'h0000FFBE3C7FE00000000003F80018041FFFFFFFFFFFFFFFFFFFFFFFFE07002F;
defparam dpb_inst_1.INIT_RAM_27 = 256'h0000FFBE3C7FE00000000003F807F8041FFFFFFFFFFFFC000003FFFFFE01002F;
defparam dpb_inst_1.INIT_RAM_28 = 256'h0000FFBE3C7FE00000000C0FF83FF8041FFFFFFFFFFFFC000003FFFFFE010C2F;
defparam dpb_inst_1.INIT_RAM_29 = 256'h0000FFBE3C7FE00000000000F83FF8041FFFFFFFFFFFFFFFFFFFFFFFFE010E2F;
defparam dpb_inst_1.INIT_RAM_2A = 256'h0000FFBE3C7FE00001800000F80018040FFFFFFFFFFFFF81F80FFFFFFE010FEF;
defparam dpb_inst_1.INIT_RAM_2B = 256'h0000FFBE387FE04000000C09F80018040FFFFFFFFFFFFC20F043FFFFFC010FEF;
defparam dpb_inst_1.INIT_RAM_2C = 256'h0000FFBE307FE00000000001F9FFF8000FFFFFFFFFFFF847FF21FFFFFC010FEF;
defparam dpb_inst_1.INIT_RAM_2D = 256'h0000FFBE287FE04000800001F800180003FFFFFFFFFFFC01FC21FFFFFC010FEF;
defparam dpb_inst_1.INIT_RAM_2E = 256'h0000FFBE387FE04000FF0C09F800180003FFFFFFFFFFFE1C0187FFFFFC010FEF;
defparam dpb_inst_1.INIT_RAM_2F = 256'h0000FFBE307FE04001FF001FF800180001FFFFFFFFFFFFF0007FFFFFF0010FEF;
defparam dpb_inst_1.INIT_RAM_30 = 256'h0000FFBE3C7FF04001FF0000FBFFF80200FFFFFFFFFFFFFFFFFFFFFFE0014FEF;
defparam dpb_inst_1.INIT_RAM_31 = 256'h0000FFBE387FF04001FF0000FBFFF802000FFFFFFFFFFFFFFFFFFFFF80014FEF;
defparam dpb_inst_1.INIT_RAM_32 = 256'h0000FFBE307FE04000FF0010FBFFF80000000000FFFFFFFFFFFC000000014FEF;
defparam dpb_inst_1.INIT_RAM_33 = 256'h0000FFBE307FF04000000000FBFFF80000000000000000000000000000014FEF;
defparam dpb_inst_1.INIT_RAM_34 = 256'h0000FFBE387FF04000040000FBFFF80000000000000000000000000000010FEF;
defparam dpb_inst_1.INIT_RAM_35 = 256'h0000FFBE307FF040000400C0FBFFF80000000000000000000000000000010FEF;
defparam dpb_inst_1.INIT_RAM_36 = 256'h0000FFBE207FF04020033800FBC2780000000000007FFFFFFFFE000000010FEF;
defparam dpb_inst_1.INIT_RAM_37 = 256'h0000FFBE207FF04000000000FBD7F800000000000040003F8103080000010FEF;
defparam dpb_inst_1.INIT_RAM_38 = 256'h0000FFBE307FF04000004000FBFFF800000000000040001F8183000000010BEF;
defparam dpb_inst_1.INIT_RAM_39 = 256'h0000FFBE207FF04000000000FB81F800000000000040881D8081000200018BEF;
defparam dpb_inst_1.INIT_RAM_3A = 256'h0000FFBE287FF0000000C0E0FBC5F800000000000040881F8081000181018FEF;
defparam dpb_inst_1.INIT_RAM_3B = 256'h0000FFBE307FF0000C000000FBFFF800000000000040001D8081000000018FEF;
defparam dpb_inst_1.INIT_RAM_3C = 256'h0000FFBE007FF00000000000FBFFF800000000000040001F8081000000018FEF;
defparam dpb_inst_1.INIT_RAM_3D = 256'h0000FFBC207FF0000000C1E0FBFFF800000000000060003F8003000000010FEF;
defparam dpb_inst_1.INIT_RAM_3E = 256'h0000FFB2207FF00000000000FBFFF80000000000000000000000000000010FF3;
defparam dpb_inst_1.INIT_RAM_3F = 256'h0000FFB2007FF00000000000FBFFF8000000000000000000000000000001B833;

DPB dpb_inst_2 (
    .DOA({dpb_inst_2_douta_w[14:0],dpb_inst_2_douta[2]}),
    .DOB({dpb_inst_2_doutb_w[14:0],dpb_inst_2_doutb[2]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[2]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[2]})
);

defparam dpb_inst_2.READ_MODE0 = 1'b1;
defparam dpb_inst_2.READ_MODE1 = 1'b1;
defparam dpb_inst_2.WRITE_MODE0 = 2'b00;
defparam dpb_inst_2.WRITE_MODE1 = 2'b00;
defparam dpb_inst_2.BIT_WIDTH_0 = 1;
defparam dpb_inst_2.BIT_WIDTH_1 = 1;
defparam dpb_inst_2.BLK_SEL_0 = 3'b000;
defparam dpb_inst_2.BLK_SEL_1 = 3'b000;
defparam dpb_inst_2.RESET_MODE = "SYNC";
defparam dpb_inst_2.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_01 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_03 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_05 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_06 = 256'h0000FF8E203FF87FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_07 = 256'h0000FFBF303FFFFF81FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_08 = 256'h0000FFBF003FFFFFFFFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_09 = 256'h0000FFBF387FF0007FFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_0A = 256'h0000FFBF307FE0000000FFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_0B = 256'h0000FFBF307FE08000000001FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_0C = 256'h0000FFBF387FE08000000000FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_0D = 256'h0000FFBF3C7FF08000000000FBFFFFFFFFFFFFFFFFFFFFFC0000000000007FFF;
defparam dpb_inst_2.INIT_RAM_0E = 256'h0000FFBF3C7FE08000300000FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FF;
defparam dpb_inst_2.INIT_RAM_0F = 256'h0000FFBF3C7FE08001000000FBFFFF8000000000000000000000000000000F1F;
defparam dpb_inst_2.INIT_RAM_10 = 256'h0000FFBF3C7FE08000000018FBFFF8000000000000000000000000000008001F;
defparam dpb_inst_2.INIT_RAM_11 = 256'h0000FFBF3C7FE08000000800FBFFF0000000000000000000000000000008001F;
defparam dpb_inst_2.INIT_RAM_12 = 256'h0000FFBF3C7FE08004000000FBFFF0060000000000000000000000000008001F;
defparam dpb_inst_2.INIT_RAM_13 = 256'h0000FFBF3C7FE08000000018FBFFF0007000FFFFFFFFFFFFFFFFFFFE0008004F;
defparam dpb_inst_2.INIT_RAM_14 = 256'h0000FFBF3C7FE08000000C00FBFFF000183FFFFFFFFFFFFFFFFFFFFFE008004F;
defparam dpb_inst_2.INIT_RAM_15 = 256'h0000FFBF387FE08000000000FBFFF00001FFFFFFFFFFFFFFFFFFFFFFF008004F;
defparam dpb_inst_2.INIT_RAM_16 = 256'h0000FFBF387FE08000000000F804700001FFFFFFFFFFFFFFFF03FFFFF008004F;
defparam dpb_inst_2.INIT_RAM_17 = 256'h0000FFBF3C7FE08000004C00F83FF00003FFFFFFFFFFFC000023FFFFFC08000F;
defparam dpb_inst_2.INIT_RAM_18 = 256'h0000FFBF387FE08002080000FBFFF00003FFFFFFFFFFFC000023FFFFFC08000F;
defparam dpb_inst_2.INIT_RAM_19 = 256'h0000FFBF3C7FE08004006000F80030000FFFFFFFFFFFFFFFFF23FFFFFE08000F;
defparam dpb_inst_2.INIT_RAM_1A = 256'h0000FFBE3C7FE08000100000F80030000FFFFFFFFFFFFFFFFFFFFFFFFE08000F;
defparam dpb_inst_2.INIT_RAM_1B = 256'h0000FFBE3C7FE08000000000F84470000FFFFFFFFFFFFC155543FFFFFE08000F;
defparam dpb_inst_2.INIT_RAM_1C = 256'h0000FFBE3C7FE08000000000FBFFF0000FFFFFFFFFFFFC000023FFFFFE08000F;
defparam dpb_inst_2.INIT_RAM_1D = 256'h0000FFBE387FE08000040000F80030001FFFFFFFFFFFFC030C23FFFFFE04000F;
defparam dpb_inst_2.INIT_RAM_1E = 256'h0000FFBE3C7FE08000000038F80010001FFFFFFFFFFFFC001C07FFFFFE04000F;
defparam dpb_inst_2.INIT_RAM_1F = 256'h0000FFBE3C7FE08000000003F8FFF0001FFFFFFFFFFFFCFFFFFFFFFFFE04000F;
defparam dpb_inst_2.INIT_RAM_20 = 256'h0000FFBE387FE08000040006F801F0001FFFFFFFFFFFFC07E003FFFFFE04002F;
defparam dpb_inst_2.INIT_RAM_21 = 256'h0000FFBE3C7FE0800000001EF80030001FFFFFFFFFFFF8460821FFFFFF04002F;
defparam dpb_inst_2.INIT_RAM_22 = 256'h0000FFBE3C7FE00000000002F80010001FFFFFFFFFFFFC218701FFFFFF04002F;
defparam dpb_inst_2.INIT_RAM_23 = 256'h0000FFBE3C7FE08000000006F80038001FFFFFFFFFFFFF803FFFFFFFFF04002F;
defparam dpb_inst_2.INIT_RAM_24 = 256'h0000FFBE3C7FE0000100003EF9FFF8001FFFFFFFFFFFFFFE07FFFFFFFF07002F;
defparam dpb_inst_2.INIT_RAM_25 = 256'h0000FFBE3C7FE0000000000FF80078001FFFFFFFFFFFFFFE27FFFFFFFF07002F;
defparam dpb_inst_2.INIT_RAM_26 = 256'h0000FFBE3C7FE00000040003F80018001FFFFFFFFFFFFFFE07FFFFFFFF07002F;
defparam dpb_inst_2.INIT_RAM_27 = 256'h0000FFBE3C7FE00000000003F80018041FFFFFFFFFFFFC000003FFFFFE01002F;
defparam dpb_inst_2.INIT_RAM_28 = 256'h0000FFBE3C7FE00000000C0FF83FF8041FFFFFFFFFFFFC000003FFFFFE010C2F;
defparam dpb_inst_2.INIT_RAM_29 = 256'h0000FFBE3C7FE00000000000F83FF8041FFFFFFFFFFFFFFFFFFFFFFFFE010E2F;
defparam dpb_inst_2.INIT_RAM_2A = 256'h0000FFBE3C7FE00000000000F80018000FFFFFFFFFFFFF80501FFFFFFE010FEF;
defparam dpb_inst_2.INIT_RAM_2B = 256'h0000FFBE387FE04000001C0FF80018040FFFFFFFFFFFFC100043FFFFFC010FEF;
defparam dpb_inst_2.INIT_RAM_2C = 256'h0000FFBE387FE00000000001F80038040FFFFFFFFFFFFC43FF21FFFFFC010FEF;
defparam dpb_inst_2.INIT_RAM_2D = 256'h0000FFBE387FE04000004001FBFFF80007FFFFFFFFFFFC43FC21FFFFFC010FEF;
defparam dpb_inst_2.INIT_RAM_2E = 256'h0000FFBE387FE040007F0C09F800180003FFFFFFFFFFFE1C0187FFFFFC010FEF;
defparam dpb_inst_2.INIT_RAM_2F = 256'h0000FFBE307FE04001FF0005F800180001FFFFFFFFFFFFF0003FFFFFF0010FEF;
defparam dpb_inst_2.INIT_RAM_30 = 256'h0000FFBE3C7FE040003F0000FBFFF80001FFFFFFFFFFFFFFFFFFFFFFE0014FEF;
defparam dpb_inst_2.INIT_RAM_31 = 256'h0000FFBE007FF04001FF0800FBFFF802001FFFFFFFFFFFFFFFFFFFFFC0014FEF;
defparam dpb_inst_2.INIT_RAM_32 = 256'h0000FFBE387FE04000FF0010FBFFF800000003FFFFFFFFFFFFFFFF0000014FEF;
defparam dpb_inst_2.INIT_RAM_33 = 256'h0000FFBE307FF04000000000FBFFF80000000000000000000000000000014FEF;
defparam dpb_inst_2.INIT_RAM_34 = 256'h0000FFBE307FF04000040000FBFFF80000000000000000000000000000010FEF;
defparam dpb_inst_2.INIT_RAM_35 = 256'h0000FFBE307FF04000040040FBFFF80000000000000000000000000000010FEF;
defparam dpb_inst_2.INIT_RAM_36 = 256'h0000FFBE207FF04000003800FB80F80000000000000000000000000000010FEF;
defparam dpb_inst_2.INIT_RAM_37 = 256'h0000FFBE207FF04000003800FBC3F800000000000040003F8003080000010FEF;
defparam dpb_inst_2.INIT_RAM_38 = 256'h0000FFBE307FF04000004000FBFFF800000000000040001F8183000000010BEF;
defparam dpb_inst_2.INIT_RAM_39 = 256'h0000FFBE207FF04000000000FB81F800000000000040801D8081000000018BEF;
defparam dpb_inst_2.INIT_RAM_3A = 256'h0000FFBE207FF00000000060FBC1F800000000000040081F8001000081018FEF;
defparam dpb_inst_2.INIT_RAM_3B = 256'h0000FFBE307FF0001C000000FBFFF800000000000040081D8081000000018FEF;
defparam dpb_inst_2.INIT_RAM_3C = 256'h0000FFBE007FF00000000000FBFFF800000000000040001F8081000000018FEF;
defparam dpb_inst_2.INIT_RAM_3D = 256'h0000FFBC207FF0000000C1E0FBFFF800000000000060003F8003000000010FEF;
defparam dpb_inst_2.INIT_RAM_3E = 256'h0000FFB2007FF00000000000FBFFF80000000000000000000000000000010FF3;
defparam dpb_inst_2.INIT_RAM_3F = 256'h0000FFB2007FF00000000000FBFFF80000000000000000000000000000018C33;

DPB dpb_inst_3 (
    .DOA({dpb_inst_3_douta_w[14:0],dpb_inst_3_douta[3]}),
    .DOB({dpb_inst_3_doutb_w[14:0],dpb_inst_3_doutb[3]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[3]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[3]})
);

defparam dpb_inst_3.READ_MODE0 = 1'b1;
defparam dpb_inst_3.READ_MODE1 = 1'b1;
defparam dpb_inst_3.WRITE_MODE0 = 2'b00;
defparam dpb_inst_3.WRITE_MODE1 = 2'b00;
defparam dpb_inst_3.BIT_WIDTH_0 = 1;
defparam dpb_inst_3.BIT_WIDTH_1 = 1;
defparam dpb_inst_3.BLK_SEL_0 = 3'b000;
defparam dpb_inst_3.BLK_SEL_1 = 3'b000;
defparam dpb_inst_3.RESET_MODE = "SYNC";
defparam dpb_inst_3.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_01 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_03 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_05 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_06 = 256'h0000FF80087FE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_07 = 256'h0000FFBF303FFFFF87FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_08 = 256'h0000FFBF003FFFFFFFFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_09 = 256'h0000FFBF387FF8007FFFFFC0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_0A = 256'h0000FFBF307FE0000007FFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_0B = 256'h0000FFBF387FE00000000003FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_0C = 256'h0000FFBF387FE08000000000FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_0D = 256'h0000FFBF3C7FF08000000000FBFFFFFFFFFFFFFFFFFFFFFC0000000000007FFF;
defparam dpb_inst_3.INIT_RAM_0E = 256'h0000FFBF3C7FE08000000000FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1FF;
defparam dpb_inst_3.INIT_RAM_0F = 256'h0000FFBF3C7FE08000040000FBFFFFFFF8000000000000000000000000000FDF;
defparam dpb_inst_3.INIT_RAM_10 = 256'h0000FFBF3C7FE08001000000FBFFF8000000000000000000000000000000001F;
defparam dpb_inst_3.INIT_RAM_11 = 256'h0000FFBF3C7FE08000000000FBFFF0000000000000000000000000000008001F;
defparam dpb_inst_3.INIT_RAM_12 = 256'h0000FFBF3C7FE08004000000FBFFF0060000000000000000000000000008001F;
defparam dpb_inst_3.INIT_RAM_13 = 256'h0000FFBF3C7FE08000000018FBFFF00060009FFFFFFFFFFFFFFFFFFA0008004F;
defparam dpb_inst_3.INIT_RAM_14 = 256'h0000FFBF387FE08000000C00FBFFF0001E1FFFFFFFFFFFFFFFFFFFFFE008004F;
defparam dpb_inst_3.INIT_RAM_15 = 256'h0000FFBF387FE08000100000FBFFF00000FFFFFFFFFFFFFFFFFFFFFFF008004F;
defparam dpb_inst_3.INIT_RAM_16 = 256'h0000FFBF387FE08000000018F800300001FFFFFFFFFFFFFFFF03FFFFF008004F;
defparam dpb_inst_3.INIT_RAM_17 = 256'h0000FFBF3C7FE08000004C00F83FF00003FFFFFFFFFFFC000023FFFFFC08000F;
defparam dpb_inst_3.INIT_RAM_18 = 256'h0000FFBF3C7FE08002000000F9FFF00003FFFFFFFFFFFC000023FFFFFC08000F;
defparam dpb_inst_3.INIT_RAM_19 = 256'h0000FFBE3C7FE08001000008F800300003FFFFFFFFFFFFFFFF23FFFFFC08000F;
defparam dpb_inst_3.INIT_RAM_1A = 256'h0000FFBE3C7FE08000000C00F80010000FFFFFFFFFFFFFFFFFFFFFFFFE08000F;
defparam dpb_inst_3.INIT_RAM_1B = 256'h0000FFBE3C7FE08000000000F80030000FFFFFFFFFFFFC000003FFFFFE08000F;
defparam dpb_inst_3.INIT_RAM_1C = 256'h0000FFBE3C7FE08000000000F9FFF0000FFFFFFFFFFFFC000023FFFFFE08000F;
defparam dpb_inst_3.INIT_RAM_1D = 256'h0000FFBE387FE08000000000F80070001FFFFFFFFFFFFE010E23FFFFFE04000F;
defparam dpb_inst_3.INIT_RAM_1E = 256'h0000FFBE387FE08000000000F80010001FFFFFFFFFFFFC403787FFFFFE04000F;
defparam dpb_inst_3.INIT_RAM_1F = 256'h0000FFBE387FE08000000000F80010001FFFFFFFFFFFFC7F80FFFFFFFE04000F;
defparam dpb_inst_3.INIT_RAM_20 = 256'h0000FFBE387FE0800004000EFBFFF0001FFFFFFFFFFFFC03E007FFFFFE04002F;
defparam dpb_inst_3.INIT_RAM_21 = 256'h0000FFBE3C7FE0800000001EF80070001FFFFFFFFFFFF8460821FFFFFF04002F;
defparam dpb_inst_3.INIT_RAM_22 = 256'h0000FFBE3C7FE00000000000F80010001FFFFFFFFFFFFC008301FFFFFF04002F;
defparam dpb_inst_3.INIT_RAM_23 = 256'h0000FFBE3C7FE0000000000EF80018001FFFFFFFFFFFFE001FFFFFFFFF04002F;
defparam dpb_inst_3.INIT_RAM_24 = 256'h0000FFBE3C7FE0800000003EF80038001FFFFFFFFFFFFFFE07FFFFFFFF04002F;
defparam dpb_inst_3.INIT_RAM_25 = 256'h0000FFBE3C7FE0000000000FFBFFF8001FFFFFFFFFFFFFFE27FFFFFFFF07002F;
defparam dpb_inst_3.INIT_RAM_26 = 256'h0000FFBE3C7FE00000040007F80018001FFFFFFFFFFFFFFE07FFFFFFFF03002F;
defparam dpb_inst_3.INIT_RAM_27 = 256'h0000FFBE3C7FE00000000007F80018041FFFFFFFFFFFFC000003FFFFFE01002F;
defparam dpb_inst_3.INIT_RAM_28 = 256'h0000FFBE3C7FE0000000000FF80018041FFFFFFFFFFFFC000003FFFFFE010C2F;
defparam dpb_inst_3.INIT_RAM_29 = 256'h0000FFBE307FE04000000003F8FFF8041FFFFFFFFFFFFFFFFFFFFFFFFE010C2F;
defparam dpb_inst_3.INIT_RAM_2A = 256'h0000FFBE3C7FE04000000001F801F8000FFFFFFFFFFFFFC0003FFFFFFE010F2F;
defparam dpb_inst_3.INIT_RAM_2B = 256'h0000FFBE387FE00000000C0FF80018040FFFFFFFFFFFFC100043FFFFFC010FEF;
defparam dpb_inst_3.INIT_RAM_2C = 256'h0000FFBE387FE00000000001F80038040FFFFFFFFFFFFC43FE21FFFFFC010FEF;
defparam dpb_inst_3.INIT_RAM_2D = 256'h0000FFBE307FE00000000001F80038000FFFFFFFFFFFFC43FC20FFFFFC010FEF;
defparam dpb_inst_3.INIT_RAM_2E = 256'h0000FFBE387FE040003F8C09FBFFF80003FFFFFFFFFFFE100083FFFFFC010FEF;
defparam dpb_inst_3.INIT_RAM_2F = 256'h0000FFBE387FE04003FF0000F800180001FFFFFFFFFFFFE0003FFFFFF0010FEF;
defparam dpb_inst_3.INIT_RAM_30 = 256'h0000FFBE3C7FE040007F0000FBFFF80001FFFFFFFFFFFFFFFFFFFFFFE0014FEF;
defparam dpb_inst_3.INIT_RAM_31 = 256'h0000FFBE007FE04001FF0800FBFFF802003FFFFFFFFFFFFFFFFFFFFFC0014FEF;
defparam dpb_inst_3.INIT_RAM_32 = 256'h0000FFBE387FF04001FF0010FBFFF80000003FFFFFFFFFFFFFFFFFF800010FEF;
defparam dpb_inst_3.INIT_RAM_33 = 256'h0000FFBE387FF04001E00000FBFFF80000000000000000000000000000014FEF;
defparam dpb_inst_3.INIT_RAM_34 = 256'h0000FFBE347FF04000000800FBFFF80000000000000000000000000000010FEF;
defparam dpb_inst_3.INIT_RAM_35 = 256'h0000FFBE307FF04000040040FBFFF80000000000000000000000000000010FEF;
defparam dpb_inst_3.INIT_RAM_36 = 256'h0000FFBE207FF04000000000FB80F80000000000000000000000000000010FEF;
defparam dpb_inst_3.INIT_RAM_37 = 256'h0000FFBE207FF04000000600FB81F800000000000040003F8003080000010BEF;
defparam dpb_inst_3.INIT_RAM_38 = 256'h0000FFBE207FF04000004040FBFFF800000000000040003F8183000000018BEF;
defparam dpb_inst_3.INIT_RAM_39 = 256'h0000FFBE207FF04000000000FBC3F800000000000040801D8081000000018BEF;
defparam dpb_inst_3.INIT_RAM_3A = 256'h0000FFBE207FF00000000060FBC1F800000000000040081F8001000081018FEF;
defparam dpb_inst_3.INIT_RAM_3B = 256'h0000FFBE307FF0001C000000FBFFF800000000000040001D8081000000018FEF;
defparam dpb_inst_3.INIT_RAM_3C = 256'h0000FFBE207FF00000000000FBFFF800000000000040001F8081000000018FEF;
defparam dpb_inst_3.INIT_RAM_3D = 256'h0000FFBC007FF000000041E0FBFFF800000000000040001F8001000000010FEF;
defparam dpb_inst_3.INIT_RAM_3E = 256'h0000FFB2007FF00000000000FBFFF80000000000000000000000000000010FF3;
defparam dpb_inst_3.INIT_RAM_3F = 256'h0000FFB2007FF00000000000FBFFF80000000000000000000000000000018C33;

DPB dpb_inst_4 (
    .DOA({dpb_inst_4_douta_w[11:0],dpb_inst_4_douta[3:0]}),
    .DOB({dpb_inst_4_doutb_w[11:0],dpb_inst_4_doutb[3:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[14],ada[13],ada[12]}),
    .BLKSELB({adb[14],adb[13],adb[12]}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[3:0]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[3:0]})
);

defparam dpb_inst_4.READ_MODE0 = 1'b1;
defparam dpb_inst_4.READ_MODE1 = 1'b1;
defparam dpb_inst_4.WRITE_MODE0 = 2'b00;
defparam dpb_inst_4.WRITE_MODE1 = 2'b00;
defparam dpb_inst_4.BIT_WIDTH_0 = 4;
defparam dpb_inst_4.BIT_WIDTH_1 = 4;
defparam dpb_inst_4.BLK_SEL_0 = 3'b100;
defparam dpb_inst_4.BLK_SEL_1 = 3'b100;
defparam dpb_inst_4.RESET_MODE = "SYNC";
defparam dpb_inst_4.INIT_RAM_00 = 256'h00000000000000000000000000000000000000000000000000000037FFFF00FF;
defparam dpb_inst_4.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_4.INIT_RAM_02 = 256'hFFFFFF00000300007F00000FFFC00000FFFFF0FFFFFFFFFFFFFFFF3300000000;
defparam dpb_inst_4.INIT_RAM_03 = 256'h0000000000000000FFFFFFFFF0FCE77000F0000000DFFFFFFFFF0000000000FF;
defparam dpb_inst_4.INIT_RAM_04 = 256'h13131313131313131313131313131313131313131313777777FFFFFE8817FFFF;
defparam dpb_inst_4.INIT_RAM_05 = 256'h7777777777777777777777777777777777313113131313131313131313131313;
defparam dpb_inst_4.INIT_RAM_06 = 256'hFFFFFF00000000000000000000000000FFFFF0FFFFFFFFFFFFFFFFFFFF777777;
defparam dpb_inst_4.INIT_RAM_07 = 256'h0000000000000000FFFFFFFFF0FE44000040000001FFFFFFFFFF0000F00000FF;
defparam dpb_inst_4.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8017FFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_09 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEFEEEEFEEFEEEEFEFEEFFF;
defparam dpb_inst_4.INIT_RAM_0A = 256'h88800000000000000000000000000000FFFFF0EEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_4.INIT_RAM_0B = 256'h0000000000000000FFFFFFFFF0F801100000000009FFFFFFFFFF0000F0000088;
defparam dpb_inst_4.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_0E = 256'h00000000000000000000000000000003FFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_0F = 256'h0000000000000000FFFFFFFFF0FC00000000000000FFFFFFFFFF000000000000;
defparam dpb_inst_4.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_12 = 256'h0000000000000000001013333FFFFFFFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_13 = 256'h0000000000000000FFFFFFFFF0F000000000000000FFFFFFFFFF000000000000;
defparam dpb_inst_4.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_16 = 256'h0333337F7FFFFFFFFFFFFFFFFFFFFFFFFFECC3FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_17 = 256'h0000000000000000FFFFFFFFF07000000000000000FFFFFFFFFF300000000000;
defparam dpb_inst_4.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFECC8991377FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_1B = 256'h0000000000000000FFFFFFFFF00000000000000000FFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_1E = 256'hFEEEC9993777FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_1F = 256'h0000000000000000FFFFFFFFF00000000000000000FFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_23 = 256'h0000000000000000FFFFFFFFF11111111000000000FFFFFEEEE88993337FFFFF;
defparam dpb_inst_4.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_27 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_2B = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_2F = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_33 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_37 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_3B = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_3F = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DPB dpb_inst_5 (
    .DOA({dpb_inst_5_douta_w[14:0],dpb_inst_5_douta[4]}),
    .DOB({dpb_inst_5_doutb_w[14:0],dpb_inst_5_doutb[4]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[4]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[4]})
);

defparam dpb_inst_5.READ_MODE0 = 1'b1;
defparam dpb_inst_5.READ_MODE1 = 1'b1;
defparam dpb_inst_5.WRITE_MODE0 = 2'b00;
defparam dpb_inst_5.WRITE_MODE1 = 2'b00;
defparam dpb_inst_5.BIT_WIDTH_0 = 1;
defparam dpb_inst_5.BIT_WIDTH_1 = 1;
defparam dpb_inst_5.BLK_SEL_0 = 3'b000;
defparam dpb_inst_5.BLK_SEL_1 = 3'b000;
defparam dpb_inst_5.RESET_MODE = "SYNC";
defparam dpb_inst_5.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_01 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_03 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_05 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_06 = 256'h0000FF80003F07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_07 = 256'h0000FFBF303FFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_08 = 256'h0000FFBF003FFFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_09 = 256'h0000FFBF387FF803FFFFFFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_0A = 256'h0000FFBF307FE0000007FFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_0B = 256'h0000FFBF307FE00000000007FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_0C = 256'h0000FFBF387FF08000000000FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_0D = 256'h0000FFBF387FE08000000000FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFF;
defparam dpb_inst_5.INIT_RAM_0E = 256'h0000FFBF387FE08000000000FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3FF;
defparam dpb_inst_5.INIT_RAM_0F = 256'h0000FFBF3C7FE08000040000FBFFFFFFFC000000000000000000000000001FDF;
defparam dpb_inst_5.INIT_RAM_10 = 256'h0000FFBF3C7FE08000000000FBFFF8000000000000000000000000000000001F;
defparam dpb_inst_5.INIT_RAM_11 = 256'h0000FFBF387FE08000000000FBFFF0000000000000000000000000000008001F;
defparam dpb_inst_5.INIT_RAM_12 = 256'h0000FFBF3C7FE08000040000FBFFF0040000000000000000000000000008001F;
defparam dpb_inst_5.INIT_RAM_13 = 256'h0000FFBF3C7FE08001000038FBFFF000600007FFFFFFFFFFFFFFFFF80008004F;
defparam dpb_inst_5.INIT_RAM_14 = 256'h0000FFBF387FE08000000C00FBFFF0001E1FFFFFFFFFFFFFFFFFFFFFE008004F;
defparam dpb_inst_5.INIT_RAM_15 = 256'h0000FFBF387FE08000000000FBFFF00000FFFFFFFFFFFFFFFFFFFFFFF008004F;
defparam dpb_inst_5.INIT_RAM_16 = 256'h0000FFBF387FE08005000038F801F00001FFFFFFFFFFFFFFFF03FFFFF008004F;
defparam dpb_inst_5.INIT_RAM_17 = 256'h0000FFBF3C7FE08000100C00F800300003FFFFFFFFFFFC000023FFFFFC08000F;
defparam dpb_inst_5.INIT_RAM_18 = 256'h0000FFBF3C7FE08006000000F8FFF00003FFFFFFFFFFFC7FFFE3FFFFFC08000F;
defparam dpb_inst_5.INIT_RAM_19 = 256'h0000FFBE3C7FE08001000008F800700003FFFFFFFFFFFFFFFF23FFFFFC08000F;
defparam dpb_inst_5.INIT_RAM_1A = 256'h0000FFBE3C7FE08000000C00F80010000FFFFFFFFFFFFFFFFF57FFFFFE0C000F;
defparam dpb_inst_5.INIT_RAM_1B = 256'h0000FFBE3C7FE08000000000F80010000FFFFFFFFFFFFC000003FFFFFE08000F;
defparam dpb_inst_5.INIT_RAM_1C = 256'h0000FFBE3C7FE08001000000F80030000FFFFFFFFFFFFC000023FFFFFE08000F;
defparam dpb_inst_5.INIT_RAM_1D = 256'h0000FFBE387FE08000000400FBFFF0001FFFFFFFFFFFFE011F23FFFFFE0C000F;
defparam dpb_inst_5.INIT_RAM_1E = 256'h0000FFBE387FE08000000000F80010001FFFFFFFFFFFFC403387FFFFFE04000F;
defparam dpb_inst_5.INIT_RAM_1F = 256'h0000FFBE3C7FE08000000000F80010001FFFFFFFFFFFFC3F807FFFFFFE04000F;
defparam dpb_inst_5.INIT_RAM_20 = 256'h0000FFBE3C7FE0800000040FF80010001FFFFFFFFFFFFC03F00FFFFFFE04002F;
defparam dpb_inst_5.INIT_RAM_21 = 256'h0000FFBE3C7FE08000000002FBFFF0001FFFFFFFFFFFF8470463FFFFFE04002F;
defparam dpb_inst_5.INIT_RAM_22 = 256'h0000FFBE387FE00000000000F80030001FFFFFFFFFFFFC008121FFFFFF04002F;
defparam dpb_inst_5.INIT_RAM_23 = 256'h0000FFBE3C7FE0000000000EF80018001FFFFFFFFFFFFE001FFFFFFFFF04002F;
defparam dpb_inst_5.INIT_RAM_24 = 256'h0000FFBE3C7FE00000000016F80030001FFFFFFFFFFFFFFE07FFFFFFFF04002F;
defparam dpb_inst_5.INIT_RAM_25 = 256'h0000FFBE3C7FE00001000003F80038001FFFFFFFFFFFFFFE27FFFFFFFF07002F;
defparam dpb_inst_5.INIT_RAM_26 = 256'h0000FFBE3C7FE0000004000FFBFFF8001FFFFFFFFFFFFFFE07FFFFFFFF01002F;
defparam dpb_inst_5.INIT_RAM_27 = 256'h0000FFBE3C7FE0000000003FF80018041FFFFFFFFFFFFC000003FFFFFE01002F;
defparam dpb_inst_5.INIT_RAM_28 = 256'h0000FFBE3C7FE00000000007F80018041FFFFFFFFFFFFC000003FFFFFE010C2F;
defparam dpb_inst_5.INIT_RAM_29 = 256'h0000FFBE307FE00000000007F84038041FFFFFFFFFFFFFFFFFFFFFFFFE010C2F;
defparam dpb_inst_5.INIT_RAM_2A = 256'h0000FFBE3C7FE04000000031FBFFF8000FFFFFFFFFFFFFE0007FFFFFFE010F2F;
defparam dpb_inst_5.INIT_RAM_2B = 256'h0000FFBE387FE00000000009F80038040FFFFFFFFFFFFE100087FFFFFE010FEF;
defparam dpb_inst_5.INIT_RAM_2C = 256'h0000FFBE387FE04000070001F80018040FFFFFFFFFFFFC43FC21FFFFFC010FEF;
defparam dpb_inst_5.INIT_RAM_2D = 256'h0000FFBE307FE00000000001F80038000FFFFFFFFFFFFC43FE21FFFFFC010FEF;
defparam dpb_inst_5.INIT_RAM_2E = 256'h0000FFBE387FE040007E8C08F844F80003FFFFFFFFFFFE000003FFFFFC010FEF;
defparam dpb_inst_5.INIT_RAM_2F = 256'h0000FFBE3C7FE04003FF0001FBFFF80001FFFFFFFFFFFFC0200FFFFFF0010FEF;
defparam dpb_inst_5.INIT_RAM_30 = 256'h0000FFBE387FE04000FF0000FBFFF80001FFFFFFFFFFFFFFFFFFFFFFF0010FEF;
defparam dpb_inst_5.INIT_RAM_31 = 256'h0000FFBE2C7FE04001FF0800FBFFF802007FFFFFFFFFFFFFFFFFFFFFC0014FEF;
defparam dpb_inst_5.INIT_RAM_32 = 256'h0000FFBE387FF04001FF0010FBFFF80000003FFFFFFFFFFFFFFFFFF800010FEF;
defparam dpb_inst_5.INIT_RAM_33 = 256'h0000FFBE387FF04000E00000FBFFF80000000000000000000000000000014FEF;
defparam dpb_inst_5.INIT_RAM_34 = 256'h0000FFBE3C7FF04000000800FBFFF80000000000000000000000000000010FEF;
defparam dpb_inst_5.INIT_RAM_35 = 256'h0000FFBE387FF04000040000FBFFF80000000000000000000000000000010FEF;
defparam dpb_inst_5.INIT_RAM_36 = 256'h0000FFBE387FF04000000000FB85F80000000000000000000000000000010FEF;
defparam dpb_inst_5.INIT_RAM_37 = 256'h0000FFBE207FF04000000600FB81F800000000000040003F8003080000010BEF;
defparam dpb_inst_5.INIT_RAM_38 = 256'h0000FFBE207FF04000000000FBFFF800000000000040003F8183000000010BEF;
defparam dpb_inst_5.INIT_RAM_39 = 256'h0000FFBE007FF04000000000FBFFF800000000000040881D8181000000010BEF;
defparam dpb_inst_5.INIT_RAM_3A = 256'h0000FFBE207FF04000000000FBC3F800000000000040001D8001000081010BEF;
defparam dpb_inst_5.INIT_RAM_3B = 256'h0000FFBE307FF0001C000000FBFFF800000000000040401D8081000000018FEF;
defparam dpb_inst_5.INIT_RAM_3C = 256'h0000FFBE207FF00000000000FBFFF800000000000040001F8081000000018FEF;
defparam dpb_inst_5.INIT_RAM_3D = 256'h0000FFBC007FF000000001C0FBFFF800000000000040001F8001000000010FEF;
defparam dpb_inst_5.INIT_RAM_3E = 256'h0000FFB0007FF00000300000FBFFF80000000000000000000000000000010FF3;
defparam dpb_inst_5.INIT_RAM_3F = 256'h0000FFB2207FF00000000000FBFFF80000000000000000000000000000010E33;

DPB dpb_inst_6 (
    .DOA({dpb_inst_6_douta_w[14:0],dpb_inst_6_douta[5]}),
    .DOB({dpb_inst_6_doutb_w[14:0],dpb_inst_6_doutb[5]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[5]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[5]})
);

defparam dpb_inst_6.READ_MODE0 = 1'b1;
defparam dpb_inst_6.READ_MODE1 = 1'b1;
defparam dpb_inst_6.WRITE_MODE0 = 2'b00;
defparam dpb_inst_6.WRITE_MODE1 = 2'b00;
defparam dpb_inst_6.BIT_WIDTH_0 = 1;
defparam dpb_inst_6.BIT_WIDTH_1 = 1;
defparam dpb_inst_6.BLK_SEL_0 = 3'b000;
defparam dpb_inst_6.BLK_SEL_1 = 3'b000;
defparam dpb_inst_6.RESET_MODE = "SYNC";
defparam dpb_inst_6.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_01 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_03 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_05 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_06 = 256'h0000FFFC003E1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_07 = 256'h0000FFBF303FFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_08 = 256'h0000FFBF003FFFFFFFC0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_09 = 256'h0000FFBF303FF81FFFFFFE1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_0A = 256'h0000FFBF387FF000003FFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_0B = 256'h0000FFBF307FE0000000003FFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_0C = 256'h0000FFBF387FF08000000000FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_0D = 256'h0000FFBF387FE08000000000FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFF;
defparam dpb_inst_6.INIT_RAM_0E = 256'h0000FFBF3C7FE08000008000FA01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7FF;
defparam dpb_inst_6.INIT_RAM_0F = 256'h0000FFBF3C7FE08001040000FBFFFFFFFFFFFFFF800000000000000000003F1F;
defparam dpb_inst_6.INIT_RAM_10 = 256'h0000FFBF387FE08000000000FBFFF8000000000000000000000000000000011F;
defparam dpb_inst_6.INIT_RAM_11 = 256'h0000FFBF387FE08000000000FBFFF0000000000000000000000000000008001F;
defparam dpb_inst_6.INIT_RAM_12 = 256'h0000FFBF3C7FE08000040000FBFFF0000000000000000000000000000008001F;
defparam dpb_inst_6.INIT_RAM_13 = 256'h0000FFBF3C7FE08005000000FBFFF001C000001FFFFFFFFFFFFFFF800008005F;
defparam dpb_inst_6.INIT_RAM_14 = 256'h0000FFBF3C7FE08000000000FBFFF000381FFFFFFFFFFFFFFFFFFFFFC008004F;
defparam dpb_inst_6.INIT_RAM_15 = 256'h0000FFBF387FE08000040000FBFFF00000FFFFFFFFFFFFFFFFFFFFFFF008004F;
defparam dpb_inst_6.INIT_RAM_16 = 256'h0000FFBF387FE08005000038F801F00001FFFFFFFFFFFFFFFF03FFFFF008004F;
defparam dpb_inst_6.INIT_RAM_17 = 256'h0000FFBF3C7FE08000100800F800300003FFFFFFFFFFFE000023FFFFFC08000F;
defparam dpb_inst_6.INIT_RAM_18 = 256'h0000FFBF387FE08000040000F800300003FFFFFFFFFFFC000023FFFFFC08000F;
defparam dpb_inst_6.INIT_RAM_19 = 256'h0000FFBF387FE08001000038FBFFF00003FFFFFFFFFFFC000023FFFFFC08000F;
defparam dpb_inst_6.INIT_RAM_1A = 256'h0000FFBE3C7FE08000004C00F80030000FFFFFFFFFFFFFFFFF03FFFFFE0C000F;
defparam dpb_inst_6.INIT_RAM_1B = 256'h0000FFBE3C7FE08000000000F80010000FFFFFFFFFFFFC000003FFFFFE08000F;
defparam dpb_inst_6.INIT_RAM_1C = 256'h0000FFBE3C7FE08001000000F80030000FFFFFFFFFFFFC000023FFFFFE00000F;
defparam dpb_inst_6.INIT_RAM_1D = 256'h0000FFBE387FE08000000C00F800F0001FFFFFFFFFFFFF811F23FFFFFE04000F;
defparam dpb_inst_6.INIT_RAM_1E = 256'h0000FFBE387FE08000000000FBFFF0001FFFFFFFFFFFFC608083FFFFFE04000F;
defparam dpb_inst_6.INIT_RAM_1F = 256'h0000FFBE3C7FE08001000000F80010001FFFFFFFFFFFFC0F001FFFFFFE04000F;
defparam dpb_inst_6.INIT_RAM_20 = 256'h0000FFBE3C7FE0800000040FF80010001FFFFFFFFFFFFC03F01FFFFFFE04002F;
defparam dpb_inst_6.INIT_RAM_21 = 256'h0000FFBE3C7FE08000000002F84470001FFFFFFFFFFFF8478663FFFFFE04002F;
defparam dpb_inst_6.INIT_RAM_22 = 256'h0000FFBE3C7FE08001000002FBFFF0001FFFFFFFFFFFFC402021FFFFFF04002F;
defparam dpb_inst_6.INIT_RAM_23 = 256'h0000FFBE3C7FE08000000C0EF80038001FFFFFFFFFFFFE000F03FFFFFF04002F;
defparam dpb_inst_6.INIT_RAM_24 = 256'h0000FFBE3C7FE00000000002F80010001FFFFFFFFFFFFFFF07FFFFFFFF04002F;
defparam dpb_inst_6.INIT_RAM_25 = 256'h0000FFBE3C7FE00001000003F80038001FFFFFFFFFFFFFFE27FFFFFFFF07002F;
defparam dpb_inst_6.INIT_RAM_26 = 256'h0000FFBE3C7FE0000000000FF844F8001FFFFFFFFFFFFFFE07FFFFFFFF03002F;
defparam dpb_inst_6.INIT_RAM_27 = 256'h0000FFBE3C7FE00000000013FBFFF8041FFFFFFFFFFFFFFFFFFFFFFFFE01002F;
defparam dpb_inst_6.INIT_RAM_28 = 256'h0000FFBE3C7FE00000000003F80018041FFFFFFFFFFFFC7FFFE3FFFFFE010C2F;
defparam dpb_inst_6.INIT_RAM_29 = 256'h0000FFBE387FE0000004000FF80018041FFFFFFFFFFFFFFFFFFFFFFFFE010C2F;
defparam dpb_inst_6.INIT_RAM_2A = 256'h0000FFBE3C7FE04000000031F9FFF8000FFFFFFFFFFFFFE0007FFFFFFE010F2F;
defparam dpb_inst_6.INIT_RAM_2B = 256'h0000FFBE387FE00000000001F80078040FFFFFFFFFFFFE000007FFFFFE010FEF;
defparam dpb_inst_6.INIT_RAM_2C = 256'h0000FFBE387FE04000000001F80038040FFFFFFFFFFFFC03FC23FFFFFC010FEF;
defparam dpb_inst_6.INIT_RAM_2D = 256'h0000FFBE3C7FE04000000019F80018000FFFFFFFFFFFF843FF21FFFFFC010FEF;
defparam dpb_inst_6.INIT_RAM_2E = 256'h0000FFBE387FE04000FC4C08F800380003FFFFFFFFFFFC200043FFFFFC010FEF;
defparam dpb_inst_6.INIT_RAM_2F = 256'h0000FFBE3C7FE04003FF0001F9FFF80001FFFFFFFFFFFFC0600FFFFFF8010FEF;
defparam dpb_inst_6.INIT_RAM_30 = 256'h0000FFBE287FE04000FF0000FBFFF80001FFFFFFFFFFFFFFFFFFFFFFF0030FEF;
defparam dpb_inst_6.INIT_RAM_31 = 256'h0000FFBE3C7FE040013F0800FBFFF80200FFFFFFFFFFFFFFFFFFFFFFE0014FEF;
defparam dpb_inst_6.INIT_RAM_32 = 256'h0000FFBE387FF04000FF0010FBFFF8010003FFFFFFFFFFFFFFFFFFFC00010FEF;
defparam dpb_inst_6.INIT_RAM_33 = 256'h0000FFBE387FF04000FC0010FBFFF80000000000000000000000000000014FEF;
defparam dpb_inst_6.INIT_RAM_34 = 256'h0000FFBE3C7FF04000000800FBFFF80000000000000000000000000000010FEF;
defparam dpb_inst_6.INIT_RAM_35 = 256'h0000FFBE387FF04000040000FBFFF80000000000000000000000000000010FEF;
defparam dpb_inst_6.INIT_RAM_36 = 256'h0000FFBE207FF04000000800FBC1F80000000000000000000000000000010FEF;
defparam dpb_inst_6.INIT_RAM_37 = 256'h0000FFBE207FF04000000800FBC1F800000000000040003F8003080000010FEF;
defparam dpb_inst_6.INIT_RAM_38 = 256'h0000FFBE207FF04000000000FBFFF800000000000040003F8183000000010BEF;
defparam dpb_inst_6.INIT_RAM_39 = 256'h0000FFBE007FF04000000000FBFFF800000000000040881D8181000000010BEF;
defparam dpb_inst_6.INIT_RAM_3A = 256'h0000FFBE207FF04000000000FBC3F800000000000040001D8001000081010BEF;
defparam dpb_inst_6.INIT_RAM_3B = 256'h0000FFBE287FF0001C30C000FBFFF800000000000040881D8181000000018FEF;
defparam dpb_inst_6.INIT_RAM_3C = 256'h0000FFBE207FF00000000040FBFFF800000000000040001D8081000000018FEF;
defparam dpb_inst_6.INIT_RAM_3D = 256'h0000FFBE007FF000000000C0FBFFF800000000000040001F8001000000010FEF;
defparam dpb_inst_6.INIT_RAM_3E = 256'h0000FFB8007FF00000300000FBFFF80000000000000000000000000000010FF3;
defparam dpb_inst_6.INIT_RAM_3F = 256'h0000FFB2007FF00000000000FBFFF80000000000000000000000000000010E33;

DPB dpb_inst_7 (
    .DOA({dpb_inst_7_douta_w[14:0],dpb_inst_7_douta[6]}),
    .DOB({dpb_inst_7_doutb_w[14:0],dpb_inst_7_doutb[6]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[6]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[6]})
);

defparam dpb_inst_7.READ_MODE0 = 1'b1;
defparam dpb_inst_7.READ_MODE1 = 1'b1;
defparam dpb_inst_7.WRITE_MODE0 = 2'b00;
defparam dpb_inst_7.WRITE_MODE1 = 2'b00;
defparam dpb_inst_7.BIT_WIDTH_0 = 1;
defparam dpb_inst_7.BIT_WIDTH_1 = 1;
defparam dpb_inst_7.BLK_SEL_0 = 3'b000;
defparam dpb_inst_7.BLK_SEL_1 = 3'b000;
defparam dpb_inst_7.RESET_MODE = "SYNC";
defparam dpb_inst_7.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_01 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_03 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_05 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_06 = 256'h0000FFFFFC007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_07 = 256'h0000FFBF303FFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_08 = 256'h0000FFBF303FFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_09 = 256'h0000FFBF303FFC3FFFFFFE1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_0A = 256'h0000FFBF387FF000007FFFFFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_0B = 256'h0000FFBF207FE000000001FFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_0C = 256'h0000FFBF307FE08000000000FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_0D = 256'h0000FFBF387FF08000000000FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_0E = 256'h0000FFBF3C7FE08000008000F801FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7FF;
defparam dpb_inst_7.INIT_RAM_0F = 256'h0000FFBF3E7FE08001000000FBFFFFFFFFFFFFFF800000000000000000003F1F;
defparam dpb_inst_7.INIT_RAM_10 = 256'h0000FFBF3C7FE08000000000FBFFFC000000000000000000000000000020031F;
defparam dpb_inst_7.INIT_RAM_11 = 256'h0000FFBF3C7FE08000008000FBFFF0000000000000000000000000000008001F;
defparam dpb_inst_7.INIT_RAM_12 = 256'h0000FFBF3C7FE08000040000FBFFF0000000000000000000000000000008005F;
defparam dpb_inst_7.INIT_RAM_13 = 256'h0000FFBF3C7FE08005000000FBFFF001C000001FFFFFFFFFFFFFFF800008005F;
defparam dpb_inst_7.INIT_RAM_14 = 256'h0000FFBF3C7FE08000000000FBFFF000381FFFFFFFFFFFFFFFFFFFFFC008004F;
defparam dpb_inst_7.INIT_RAM_15 = 256'h0000FFBF3C7FE08000040000FBFFF00000FFFFFFFFFFFFFFFFFFFFFFE008004F;
defparam dpb_inst_7.INIT_RAM_16 = 256'h0000FFBF387FE08005000000FBFFF00001FFFFFFFFFFFFFFFFFFFFFFF008004F;
defparam dpb_inst_7.INIT_RAM_17 = 256'h0000FFBF3C7FE08000300000F800300003FFFFFFFFFFFFFFFF23FFFFFC08000F;
defparam dpb_inst_7.INIT_RAM_18 = 256'h0000FFBF387FE08000040000F800300003FFFFFFFFFFFC000023FFFFFC08000F;
defparam dpb_inst_7.INIT_RAM_19 = 256'h0000FFBF3C7FE08001000018F800700003FFFFFFFFFFFC000023FFFFFC08000F;
defparam dpb_inst_7.INIT_RAM_1A = 256'h0000FFBE3C7FE08000000000FBFFF0000FFFFFFFFFFFFFFFFF03FFFFFE08000F;
defparam dpb_inst_7.INIT_RAM_1B = 256'h0000FFBE3C7FE08000000000F80030000FFFFFFFFFFFFC000003FFFFFE0C000F;
defparam dpb_inst_7.INIT_RAM_1C = 256'h0000FFBE3C7FE08001000018F80010000FFFFFFFFFFFFC000023FFFFFE00000F;
defparam dpb_inst_7.INIT_RAM_1D = 256'h0000FFBE387FE08000000C00F80070001FFFFFFFFFFFFF811F23FFFFFE04000F;
defparam dpb_inst_7.INIT_RAM_1E = 256'h0000FFBE387FE08000000000F847F0001FFFFFFFFFFFFC308003FFFFFE04000F;
defparam dpb_inst_7.INIT_RAM_1F = 256'h0000FFBE3C7FE08001000018FBFFF0001FFFFFFFFFFFFC06000FFFFFFE04000F;
defparam dpb_inst_7.INIT_RAM_20 = 256'h0000FFBE3C7FE08000000C0EF80010081FFFFFFFFFFFFC07FC7FFFFFFE04002F;
defparam dpb_inst_7.INIT_RAM_21 = 256'h0000FFBE3C7FE08000000002F80030001FFFFFFFFFFFFC4783C3FFFFFE04002F;
defparam dpb_inst_7.INIT_RAM_22 = 256'h0000FFBE3C7FE08001000002F9FFF0001FFFFFFFFFFFFC402021FFFFFF04002F;
defparam dpb_inst_7.INIT_RAM_23 = 256'h0000FFBE3C7FE0000000080EF80078001FFFFFFFFFFFFE000F01FFFFFF04002F;
defparam dpb_inst_7.INIT_RAM_24 = 256'h0000FFBE3C7FE00000000002F80038001FFFFFFFFFFFFFFFFFFFFFFFFF04002F;
defparam dpb_inst_7.INIT_RAM_25 = 256'h0000FFBE3C7FE00001000003F80018001FFFFFFFFFFFFFFE27FFFFFFFF07002F;
defparam dpb_inst_7.INIT_RAM_26 = 256'h0000FFBE3C7FE0000000000FF80038001FFFFFFFFFFFFFFE07FFFFFFFF07002F;
defparam dpb_inst_7.INIT_RAM_27 = 256'h0000FFBE3C7FE00000000013F9FFF8041FFFFFFFFFFFFFFFFFFFFFFFFE03002F;
defparam dpb_inst_7.INIT_RAM_28 = 256'h0000FFBE3C7FE00000000003F80018041FFFFFFFFFFFFC155543FFFFFE01082F;
defparam dpb_inst_7.INIT_RAM_29 = 256'h0000FFBE387FE0400000080FF80018041FFFFFFFFFFFFC000003FFFFFE010C2F;
defparam dpb_inst_7.INIT_RAM_2A = 256'h0000FFBE387FE04000000031F80018041FFFFFFFFFFFFFF000FFFFFFFE010F2F;
defparam dpb_inst_7.INIT_RAM_2B = 256'h0000FFBE387FE00000000001FBFFF8040FFFFFFFFFFFFE040107FFFFFE010FEF;
defparam dpb_inst_7.INIT_RAM_2C = 256'h0000FFBE387FE04000000001F80078040FFFFFFFFFFFFC03FC23FFFFFC010FEF;
defparam dpb_inst_7.INIT_RAM_2D = 256'h0000FFBE3C7FE04000000019F80018000FFFFFFFFFFFF843FF21FFFFFC010FEF;
defparam dpb_inst_7.INIT_RAM_2E = 256'h0000FFBE387FE04000F80001F800180003FFFFFFFFFFFC21F843FFFFFC010FEF;
defparam dpb_inst_7.INIT_RAM_2F = 256'h0000FFBE347FE04001FF4001F800380003FFFFFFFFFFFF83FC0FFFFFFC010FEF;
defparam dpb_inst_7.INIT_RAM_30 = 256'h0000FFBE287FE04000FF0018FBFFF80001FFFFFFFFFFFFFF9FFFFFFFF0014FEF;
defparam dpb_inst_7.INIT_RAM_31 = 256'h0000FFBE3C7FE040013F0800FBFFF80200FFFFFFFFFFFFFFFFFFFFFFE0014FEF;
defparam dpb_inst_7.INIT_RAM_32 = 256'h0000FFBE387FE04000FF0010FBFFF8000003FFFFFFFFFFFFFFFFFFFE00010FEF;
defparam dpb_inst_7.INIT_RAM_33 = 256'h0000FFBE387FF04000FF0010FBFFF8000000000000007E060000000000014FEF;
defparam dpb_inst_7.INIT_RAM_34 = 256'h0000FFBE3C7FF04000000800FBFFF80000000000000000000000000000010FEF;
defparam dpb_inst_7.INIT_RAM_35 = 256'h0000FFBE387FF04000040040FBFFF80000000000000000000000000000010FEF;
defparam dpb_inst_7.INIT_RAM_36 = 256'h0000FFBE207FF04000000800FBC1F80000000000000000000000000000010FEF;
defparam dpb_inst_7.INIT_RAM_37 = 256'h0000FFBE207FF04000000000FBC0F800000000000040003FC003080000010FEF;
defparam dpb_inst_7.INIT_RAM_38 = 256'h0000FFBE207FF04000000400FBFFF800000000000040003F81830800000103EF;
defparam dpb_inst_7.INIT_RAM_39 = 256'h0000FFBE207FF04000000000FBFFF800000000000040001F8081000000018BEF;
defparam dpb_inst_7.INIT_RAM_3A = 256'h0000FFBE207FF04000000000FBC3F800000000000040881D8181000081018BEF;
defparam dpb_inst_7.INIT_RAM_3B = 256'h0000FFBE287FF0000C30C000FBFFF800000000000040881D8181000000018FEF;
defparam dpb_inst_7.INIT_RAM_3C = 256'h0000FFBE007FF00000000040FBFFF800000000000040001D8081000000018FEF;
defparam dpb_inst_7.INIT_RAM_3D = 256'h0000FFB2007FF00000000000FBFFF800000000000040001F8081000000010FEF;
defparam dpb_inst_7.INIT_RAM_3E = 256'h0000FFBE307FF0000030C100FBFFF80000000000007FFFFFFFFF000000010FF3;
defparam dpb_inst_7.INIT_RAM_3F = 256'h0000FFB2007FF00000000040FBFFF80000000000000000000000000000018E33;

DPB dpb_inst_8 (
    .DOA({dpb_inst_8_douta_w[14:0],dpb_inst_8_douta[7]}),
    .DOB({dpb_inst_8_doutb_w[14:0],dpb_inst_8_doutb[7]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[7]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[7]})
);

defparam dpb_inst_8.READ_MODE0 = 1'b1;
defparam dpb_inst_8.READ_MODE1 = 1'b1;
defparam dpb_inst_8.WRITE_MODE0 = 2'b00;
defparam dpb_inst_8.WRITE_MODE1 = 2'b00;
defparam dpb_inst_8.BIT_WIDTH_0 = 1;
defparam dpb_inst_8.BIT_WIDTH_1 = 1;
defparam dpb_inst_8.BLK_SEL_0 = 3'b000;
defparam dpb_inst_8.BLK_SEL_1 = 3'b000;
defparam dpb_inst_8.RESET_MODE = "SYNC";
defparam dpb_inst_8.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_01 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_03 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_05 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_06 = 256'h0000FFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_07 = 256'h0000FFBE303FFF03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_08 = 256'h0000FFBF203FFFFFFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_09 = 256'h0000FFBF303FFFFFFFFFE1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_0A = 256'h0000FFBF387FF00001FFFFFF87FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_0B = 256'h0000FFBF207FE000000001FFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_0C = 256'h0000FFBF307FE08000000000FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_0D = 256'h0000FFBF387FF08000000000FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_0E = 256'h0000FFBF3C7FF08000000000F800000000000001FFFFFFFFFFFFFFFFFFFF8FFF;
defparam dpb_inst_8.INIT_RAM_0F = 256'h0000FFBF3F7FE08001000C00FBFFFFFFFFFFFFFFFFFFFFFFE000000000007E3F;
defparam dpb_inst_8.INIT_RAM_10 = 256'h0000FFBF3C7FE08000000000FBFFFE000000000000000000000000000020031F;
defparam dpb_inst_8.INIT_RAM_11 = 256'h0000FFBF3C7FE08000000000FBFFF0000000000000000000000000000008001F;
defparam dpb_inst_8.INIT_RAM_12 = 256'h0000FFBF3C7FE08000000C00FBFFF0000000000000000000000000000008001F;
defparam dpb_inst_8.INIT_RAM_13 = 256'h0000FFBF3C7FE08000000000FBFFF003C000000007FFFFFFFFFF00000008001F;
defparam dpb_inst_8.INIT_RAM_14 = 256'h0000FFBF3C7FE08000000000FBFFF000380FFFFFFFFFFFFFFFFFFFFFC008004F;
defparam dpb_inst_8.INIT_RAM_15 = 256'h0000FFBF3C7FE08000040000FBFFF00000FFFFFFFFFFFFFFFFFFFFFFE008004F;
defparam dpb_inst_8.INIT_RAM_16 = 256'h0000FFBF307FE08000000000FBFFF00001FFFFFFFFFFFFFFFFFFFFFFF008004F;
defparam dpb_inst_8.INIT_RAM_17 = 256'h0000FFBF3C7FE08000000000FBFFF00003FFFFFFFFFFFFFFFF03FFFFFC08004F;
defparam dpb_inst_8.INIT_RAM_18 = 256'h0000FFBF387FE08000040000F800300003FFFFFFFFFFFC000023FFFFFC08000F;
defparam dpb_inst_8.INIT_RAM_19 = 256'h0000FFBF3C7FE08005000018F800300003FFFFFFFFFFFC000023FFFFFC08000F;
defparam dpb_inst_8.INIT_RAM_1A = 256'h0000FFBE3C7FE08000000000F9FFF0000FFFFFFFFFFFFFFFFF03FFFFFE08000F;
defparam dpb_inst_8.INIT_RAM_1B = 256'h0000FFBE3C7FE08000000000F80070000FFFFFFFFFFFFC000003FFFFFE0C000F;
defparam dpb_inst_8.INIT_RAM_1C = 256'h0000FFBE3C7FE08000000038F80030000FFFFFFFFFFFFC3FFFE3FFFFFE08000F;
defparam dpb_inst_8.INIT_RAM_1D = 256'h0000FFBE387FE08000000000F80010001FFFFFFFFFFFFFE01F23FFFFFE04000F;
defparam dpb_inst_8.INIT_RAM_1E = 256'h0000FFBE387FE08000040000F803F0001FFFFFFFFFFFFC308043FFFFFE04000F;
defparam dpb_inst_8.INIT_RAM_1F = 256'h0000FFBE3C7FE08001000018F9FFF0001FFFFFFFFFFFFC06000FFFFFFE04000F;
defparam dpb_inst_8.INIT_RAM_20 = 256'h0000FFBE3C7FE08000000006F80010001FFFFFFFFFFFFE0FFE7FFFFFFE04002F;
defparam dpb_inst_8.INIT_RAM_21 = 256'h0000FFBE387FE08000040002F80010001FFFFFFFFFFFFC478003FFFFFE04002F;
defparam dpb_inst_8.INIT_RAM_22 = 256'h0000FFBE3C7FE08001000002F80030001FFFFFFFFFFFF8401021FFFFFF04002F;
defparam dpb_inst_8.INIT_RAM_23 = 256'h0000FFBE3C7FE0000000080FFBFFF8001FFFFFFFFFFFFC040F01FFFFFF04002F;
defparam dpb_inst_8.INIT_RAM_24 = 256'h0000FFBE3C7FE00000000002F80078001FFFFFFFFFFFFFFFFFFFFFFFFF04002F;
defparam dpb_inst_8.INIT_RAM_25 = 256'h0000FFBE3C7FE00001000003F80018001FFFFFFFFFFFFFFE27FFFFFFFF07002F;
defparam dpb_inst_8.INIT_RAM_26 = 256'h0000FFBE3C7FE00000000C0FF80018001FFFFFFFFFFFFFFE27FFFFFFFF07002F;
defparam dpb_inst_8.INIT_RAM_27 = 256'h0000FFBE3C7FE00000000003F803F8001FFFFFFFFFFFFFFFFFFFFFFFFE07002F;
defparam dpb_inst_8.INIT_RAM_28 = 256'h0000FFBE3C7FE00001800001FBFFF8041FFFFFFFFFFFFC000003FFFFFE01002F;
defparam dpb_inst_8.INIT_RAM_29 = 256'h0000FFBE387FE0000000080FF80018041FFFFFFFFFFFFC000003FFFFFE010C2F;
defparam dpb_inst_8.INIT_RAM_2A = 256'h0000FFBE387FE00000000011F80018041FFFFFFFFFFFFFF800FFFFFFFE010F2F;
defparam dpb_inst_8.INIT_RAM_2B = 256'h0000FFBE387FE04001000001F80018000FFFFFFFFFFFFF830C0FFFFFFE010FEF;
defparam dpb_inst_8.INIT_RAM_2C = 256'h0000FFBE3C7FE0400000000FFBFFF8040FFFFFFFFFFFFC21F843FFFFFC010FEF;
defparam dpb_inst_8.INIT_RAM_2D = 256'h0000FFBE387FE04000000039F80038000FFFFFFFFFFFF84FFF21FFFFFC010FEF;
defparam dpb_inst_8.INIT_RAM_2E = 256'h0000FFBE387FE04000F80001F800180003FFFFFFFFFFFC21F843FFFFFC010FEF;
defparam dpb_inst_8.INIT_RAM_2F = 256'h0000FFBE307FE04000FF4001F800380003FFFFFFFFFFFF82560FFFFFFC010FEF;
defparam dpb_inst_8.INIT_RAM_30 = 256'h0000FFBE387FE04000FF001FF800F80001FFFFFFFFFFFFFC01FFFFFFF0010FEF;
defparam dpb_inst_8.INIT_RAM_31 = 256'h0000FFBE387FE040013F0800FBFFF80200FFFFFFFFFFFFFFFFFFFFFFE0010FEF;
defparam dpb_inst_8.INIT_RAM_32 = 256'h0000FFBE387FE04001FF0010FBFFF8000007FFFFFFFFFFFFFFFFFFFE00010FEF;
defparam dpb_inst_8.INIT_RAM_33 = 256'h0000FFBE387FF04000FF0010FBFFF8000000000000007F0E0000000000014FEF;
defparam dpb_inst_8.INIT_RAM_34 = 256'h0000FFBE347FF04000000800FBFFF80000000000000000000000000000010FEF;
defparam dpb_inst_8.INIT_RAM_35 = 256'h0000FFBE387FF04000040100FBFFF80000000000000000000000000000010FEF;
defparam dpb_inst_8.INIT_RAM_36 = 256'h0000FFBE307FF04000000100FBE3F80000000000000000000000000000010FEF;
defparam dpb_inst_8.INIT_RAM_37 = 256'h0000FFBE207FF04000010400FBC2F80000000000007FFFFFFFFF080000010FEF;
defparam dpb_inst_8.INIT_RAM_38 = 256'h0000FFBE207FF04000000400FBFFF800000000000040003F81830800000103EF;
defparam dpb_inst_8.INIT_RAM_39 = 256'h0000FFBE207FF04000000000FBFFF800000000000040001D8081000000010BEF;
defparam dpb_inst_8.INIT_RAM_3A = 256'h0000FFBE007FF04000000000FB85F800000000000040881D8081000200010BEF;
defparam dpb_inst_8.INIT_RAM_3B = 256'h0000FFBE287FF0000000C1E0FBC3F800000000000040081F8001000201018FEF;
defparam dpb_inst_8.INIT_RAM_3C = 256'h0000FFBE107FF00000000040FBFFF800000000000040001F8081000000018FEF;
defparam dpb_inst_8.INIT_RAM_3D = 256'h0000FFBA007FF00000000000FBFFF800000000000040001F8081000000010FEF;
defparam dpb_inst_8.INIT_RAM_3E = 256'h0000FFBE007FF0000030C180FBFFF80000000000007FFFFFFFFF000000010FFF;
defparam dpb_inst_8.INIT_RAM_3F = 256'h0000FFB2207FF00000000040FBFFF80000000000000000000000000000018FF3;

DPB dpb_inst_9 (
    .DOA({dpb_inst_9_douta_w[11:0],dpb_inst_9_douta[7:4]}),
    .DOB({dpb_inst_9_doutb_w[11:0],dpb_inst_9_doutb[7:4]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[14],ada[13],ada[12]}),
    .BLKSELB({adb[14],adb[13],adb[12]}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[7:4]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[7:4]})
);

defparam dpb_inst_9.READ_MODE0 = 1'b1;
defparam dpb_inst_9.READ_MODE1 = 1'b1;
defparam dpb_inst_9.WRITE_MODE0 = 2'b00;
defparam dpb_inst_9.WRITE_MODE1 = 2'b00;
defparam dpb_inst_9.BIT_WIDTH_0 = 4;
defparam dpb_inst_9.BIT_WIDTH_1 = 4;
defparam dpb_inst_9.BLK_SEL_0 = 3'b100;
defparam dpb_inst_9.BLK_SEL_1 = 3'b100;
defparam dpb_inst_9.RESET_MODE = "SYNC";
defparam dpb_inst_9.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000080000007FF00FF;
defparam dpb_inst_9.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_02 = 256'h7FFF7700000000000100000017100000FFFFF0FFFFFFFFFFFFFFFF0000000000;
defparam dpb_inst_9.INIT_RAM_03 = 256'h0000000000000000FFFFFFFFF0F9CE80001000000FFFFFFFFFFF000060000037;
defparam dpb_inst_9.INIT_RAM_04 = 256'h00000000000000000000000000000000000000000000000000017FFFFFE801FF;
defparam dpb_inst_9.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_9.INIT_RAM_06 = 256'hFFFFFF00006E00008800000000000000FFFFF0FFFFFFFFFFFFFFFFFF31000000;
defparam dpb_inst_9.INIT_RAM_07 = 256'h0000000000000000FFFFFFFFF0F700000080000008FFFFFFFFFF0000300000FF;
defparam dpb_inst_9.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC033FFFFFFF;
defparam dpb_inst_9.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_0A = 256'hFFFFEE00000000000000000000000000FFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_0B = 256'h0000000000000000FFFFFFFFF0F300C0000000000FFFFFFFFFFF0000F00000FF;
defparam dpb_inst_9.INIT_RAM_0C = 256'h333333333333333333333333333333333333333333333333337FFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_0D = 256'h3333333333333333333333333333333333333333333333333333333333333333;
defparam dpb_inst_9.INIT_RAM_0E = 256'h00000000000000000000000000000000FFFFF013333333333333333333333333;
defparam dpb_inst_9.INIT_RAM_0F = 256'h0000000000000000FFFFFFFFF0FF00000000000000FFFFFFFFFF0000F0000000;
defparam dpb_inst_9.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_12 = 256'h0000000000000000000000000000113FFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_13 = 256'h0000000000000000FFFFFFFFF0F300000000000000FFFFFFFFFF000000000000;
defparam dpb_inst_9.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_16 = 256'h00000000001113777FFFFFFFFFFFFFFFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_17 = 256'h0000000000000000FFFFFFFFF0E000000000000000FFFFFFFFFF000000000000;
defparam dpb_inst_9.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFEEEC9913337FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_1B = 256'h0000000000000000FFFFFFFFF00000000000000000FFFFFFFFFFF73113373FFF;
defparam dpb_inst_9.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_1E = 256'hFFFFFFFFFEECCC93337FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_1F = 256'h0000000000000000FFFFFFFFF00000000000000000FFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_22 = 256'h3377FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_23 = 256'h0000000000000000FFFFFFFFF00000000000000000FFFFFFFFFFFFFFFFECC013;
defparam dpb_inst_9.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_27 = 256'h0000000000000000FFFFFFFFFFFFFFFFF7713113139999913777FFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_2B = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_2F = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_33 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_37 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_3B = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_3F = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ada[14]),
  .CLK(clka),
  .CE(cea_w)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(dff_q_0),
  .CLK(clka),
  .CE(ocea)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(adb[14]),
  .CLK(clkb),
  .CE(ceb_w)
);
DFFE dff_inst_3 (
  .Q(dff_q_3),
  .D(dff_q_2),
  .CLK(clkb),
  .CE(oceb)
);
MUX2 mux_inst_4 (
  .O(douta[0]),
  .I0(dpb_inst_0_douta[0]),
  .I1(dpb_inst_4_douta[0]),
  .S0(dff_q_1)
);
MUX2 mux_inst_9 (
  .O(douta[1]),
  .I0(dpb_inst_1_douta[1]),
  .I1(dpb_inst_4_douta[1]),
  .S0(dff_q_1)
);
MUX2 mux_inst_14 (
  .O(douta[2]),
  .I0(dpb_inst_2_douta[2]),
  .I1(dpb_inst_4_douta[2]),
  .S0(dff_q_1)
);
MUX2 mux_inst_19 (
  .O(douta[3]),
  .I0(dpb_inst_3_douta[3]),
  .I1(dpb_inst_4_douta[3]),
  .S0(dff_q_1)
);
MUX2 mux_inst_24 (
  .O(douta[4]),
  .I0(dpb_inst_5_douta[4]),
  .I1(dpb_inst_9_douta[4]),
  .S0(dff_q_1)
);
MUX2 mux_inst_29 (
  .O(douta[5]),
  .I0(dpb_inst_6_douta[5]),
  .I1(dpb_inst_9_douta[5]),
  .S0(dff_q_1)
);
MUX2 mux_inst_34 (
  .O(douta[6]),
  .I0(dpb_inst_7_douta[6]),
  .I1(dpb_inst_9_douta[6]),
  .S0(dff_q_1)
);
MUX2 mux_inst_39 (
  .O(douta[7]),
  .I0(dpb_inst_8_douta[7]),
  .I1(dpb_inst_9_douta[7]),
  .S0(dff_q_1)
);
MUX2 mux_inst_44 (
  .O(doutb[0]),
  .I0(dpb_inst_0_doutb[0]),
  .I1(dpb_inst_4_doutb[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_49 (
  .O(doutb[1]),
  .I0(dpb_inst_1_doutb[1]),
  .I1(dpb_inst_4_doutb[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_54 (
  .O(doutb[2]),
  .I0(dpb_inst_2_doutb[2]),
  .I1(dpb_inst_4_doutb[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_59 (
  .O(doutb[3]),
  .I0(dpb_inst_3_doutb[3]),
  .I1(dpb_inst_4_doutb[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_64 (
  .O(doutb[4]),
  .I0(dpb_inst_5_doutb[4]),
  .I1(dpb_inst_9_doutb[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_69 (
  .O(doutb[5]),
  .I0(dpb_inst_6_doutb[5]),
  .I1(dpb_inst_9_doutb[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_74 (
  .O(doutb[6]),
  .I0(dpb_inst_7_doutb[6]),
  .I1(dpb_inst_9_doutb[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_79 (
  .O(doutb[7]),
  .I0(dpb_inst_8_doutb[7]),
  .I1(dpb_inst_9_doutb[7]),
  .S0(dff_q_3)
);
endmodule //blk_mem_gen_4
