// This program was cloned from: https://github.com/sdmay24-21/ASIC-GuitarPedal
// License: Apache License 2.0

  module our;
     initial begin $display("Hello World"); $finish; end
  endmodule
