// This program was cloned from: https://github.com/Nilesh002/Multiplication-and-Accumulation-Unit-MAC-
// License: MIT License

module adder16(a,b,s);
input [15:0]a,b;
output [15:0]s;

assign s=a+b;

endmodule
