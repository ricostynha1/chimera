// This program was cloned from: https://github.com/neelkshah/MIPS-Processor
// License: GNU General Public License v3.0

module DataMemory32(clk, MemRead, ReadAddress, ReadData, MemWrite, WriteAddress, WriteData);
	input MemRead, MemWrite, clk;
	input [31:0] ReadAddress, WriteAddress;
	input [31:0] WriteData;
	output reg [31:0] ReadData;
	reg [31:0] data [0:31];
	integer raddr, waddr;
	initial
		begin
			data[0] = 32'b00000000000000000000000000000000;  
			data[1] = 32'b00000000000000000000000000000000;
			data[2] = 32'b00000000000000000000000000000000;
			data[3] = 32'b00000000000000000000000000000000;  
			data[4] = 32'b00000000000000000000000000000000;  
			data[5] = 32'b00000000000000000000000000000000;  
			data[6] = 32'b00000000000000000000000000000000;  
			data[7] = 32'b00000000000000000000000000000000;  
			data[8] = 32'b00000000000000000000000000000000;  
			data[9] = 32'b00000000000000000000000000000000;  
			data[10] = 32'b00000000000000000000000000000000;  
			data[11] = 32'b00000000000000000000000000000000;  
			data[12] = 32'b00000000000000000000000000000000;  
			data[13] = 32'b00000000000000000000000000000000;  
			data[14] = 32'b00000000000000000000000000000000;  
			data[15] = 32'b00000000000000000000000000000000;  
			data[16] = 32'b00000000000000000000000000000000;  
			data[17] = 32'b00000000000000000000000000000000;  
			data[18] = 32'b00000000000000000000000000000000;  
			data[19] = 32'b00000000000000000000000000000000;  
			data[20] = 32'b00000000000000000000000000000000;  
			data[21] = 32'b00000000000000000000000000000000;  
			data[22] = 32'b00000000000000000000000000000000;  
			data[23] = 32'b00000000000000000000000000000000;  
			data[24] = 32'b00000000000000000000000000000000;  
			data[25] = 32'b00000000000000000000000000000000;  
			data[26] = 32'b00000000000000000000000000000000;  
			data[27] = 32'b00000000000000000000000000000000;  
			data[28] = 32'b00000000000000000000000000000000;  
			data[29] = 32'b00000000000000000000000000000000;  
			data[30] = 32'b00000000000000000000000000000000;  
			data[31] = 32'b00000000000000000000000000000000;    
		end
		
	always @(posedge clk) begin
		raddr = ReadAddress;
		waddr = WriteAddress;
		if(MemRead)
			ReadData = data[raddr/4];
		else if(MemWrite)
			data[waddr/4] = WriteData;
	end
	
endmodule