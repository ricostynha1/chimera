// This program was cloned from: https://github.com/Nilesh002/Multiplication-and-Accumulation-Unit-MAC-
// License: MIT License

module add32(a,b,s);
input [31:0]a,b;
output [31:0]s;

assign s=a+b;

endmodule
