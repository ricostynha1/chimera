// This program was cloned from: https://github.com/waynezv/FPGA_Ultrasound
// License: GNU General Public License v3.0

// Jagadeesh Vasudevamurthy data_acquis_controller_X99.v
// Please do not remove the header
// Char array passed is as follows
//--------------------------------------
//0:000000 011010110111
//1:000001 010101110111
//2:000010 010001001000
//3:000011 001100110010
//4:000100 001000111011
//5:000101 000101101011
//6:000110 000011000110
//7:000111 000001010001
//8:001000 000000001111
//9:001001 000000000010
//10:001010 000000101001
//11:001011 000010000101
//12:001100 000100010010
//13:001101 000111001110
//14:001110 001010110010
//15:001111 001110111001
//16:010000 010011011101
//17:010001 011000010110
//18:010010 011101011011
//19:010011 100010100101
//20:010100 100111101010
//21:010101 101100100011
//22:010110 110001000111
//23:010111 110101001110
//24:011000 111000110010
//25:011001 111011101110
//26:011010 111101111011
//27:011011 111111010111
//28:011100 111111111110
//29:011101 111111110001
//30:011110 111110101111
//31:011111 111100111010
//32:100000 111010010101
//33:100001 110111000101
//34:100010 110011001110
//35:100011 101110111000
//36:100100 101010001001
//37:100101 100101001001
//38:100110 100000000000
// default NOT given
// Parallel mux
//--------------------------------------
// PLA starts now
module data_acquis_controller_X99(a,o);
	input[5:0]  a;
	output reg[11:0]  o;
	always @(a)
	begin
		case(a)
			6'b000000: o = 12'b011010110111;
			6'b000001: o = 12'b010101110111;
			6'b000010: o = 12'b010001001000;
			6'b000011: o = 12'b001100110010;
			6'b000100: o = 12'b001000111011;
			6'b000101: o = 12'b000101101011;
			6'b000110: o = 12'b000011000110;
			6'b000111: o = 12'b000001010001;
			6'b001000: o = 12'b000000001111;
			6'b001001: o = 12'b000000000010;
			6'b001010: o = 12'b000000101001;
			6'b001011: o = 12'b000010000101;
			6'b001100: o = 12'b000100010010;
			6'b001101: o = 12'b000111001110;
			6'b001110: o = 12'b001010110010;
			6'b001111: o = 12'b001110111001;
			6'b010000: o = 12'b010011011101;
			6'b010001: o = 12'b011000010110;
			6'b010010: o = 12'b011101011011;
			6'b010011: o = 12'b100010100101;
			6'b010100: o = 12'b100111101010;
			6'b010101: o = 12'b101100100011;
			6'b010110: o = 12'b110001000111;
			6'b010111: o = 12'b110101001110;
			6'b011000: o = 12'b111000110010;
			6'b011001: o = 12'b111011101110;
			6'b011010: o = 12'b111101111011;
			6'b011011: o = 12'b111111010111;
			6'b011100: o = 12'b111111111110;
			6'b011101: o = 12'b111111110001;
			6'b011110: o = 12'b111110101111;
			6'b011111: o = 12'b111100111010;
			6'b100000: o = 12'b111010010101;
			6'b100001: o = 12'b110111000101;
			6'b100010: o = 12'b110011001110;
			6'b100011: o = 12'b101110111000;
			6'b100100: o = 12'b101010001001;
			6'b100101: o = 12'b100101001001;
			6'b100110: o = 12'b100000000000;
// defaults of ALL_0 and ALL_X are never routine to input pla. ALL_X,ALL_1 are expanded by me. Output never has default
//			 Parallel mux
		endcase
	end
endmodule
