// This program was cloned from: https://github.com/apuder/TRS-IO
// License: GNU General Public License v3.0

//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.9 Beta-4 Education
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Device Version: C
//Created Time: Fri Feb 23 00:59:57 2024

module Gowin_DPB2 (douta, doutb, clka, ocea, cea, reseta, wrea, clkb, oceb, ceb, resetb, wreb, ada, dina, adb, dinb);

output [7:0] douta;
output [7:0] doutb;
input clka;
input ocea;
input cea;
input reseta;
input wrea;
input clkb;
input oceb;
input ceb;
input resetb;
input wreb;
input [10:0] ada;
input [7:0] dina;
input [10:0] adb;
input [7:0] dinb;

wire [7:0] dpb_inst_0_douta_w;
wire [7:0] dpb_inst_0_doutb_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

DPB dpb_inst_0 (
    .DOA({dpb_inst_0_douta_w[7:0],douta[7:0]}),
    .DOB({dpb_inst_0_doutb_w[7:0],doutb[7:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[7:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[7:0]})
);

defparam dpb_inst_0.READ_MODE0 = 1'b1;
defparam dpb_inst_0.READ_MODE1 = 1'b1;
defparam dpb_inst_0.WRITE_MODE0 = 2'b00;
defparam dpb_inst_0.WRITE_MODE1 = 2'b00;
defparam dpb_inst_0.BIT_WIDTH_0 = 8;
defparam dpb_inst_0.BIT_WIDTH_1 = 8;
defparam dpb_inst_0.BLK_SEL_0 = 3'b000;
defparam dpb_inst_0.BLK_SEL_1 = 3'b000;
defparam dpb_inst_0.RESET_MODE = "SYNC";
defparam dpb_inst_0.INIT_RAM_00 = 256'h5431FF3031335E30BF3372331B335334C2347DC9300D31F8D3ECD3003E56EDF3;
defparam dpb_inst_0.INIT_RAM_01 = 256'hFB34443029310031373C40345730873041335B32E73444301F335B000031B631;
defparam dpb_inst_0.INIT_RAM_02 = 256'h4733533061335B332B3353305D30F933723137332333533CC0345734D8347D32;
defparam dpb_inst_0.INIT_RAM_03 = 256'h1C315432D33444307F335B315431BD32DD34443079335E337231373CC0345733;
defparam dpb_inst_0.INIT_RAM_04 = 256'h78C1335631D6327834443467C9309431D90839000021EB08D93065335B306131;
defparam dpb_inst_0.INIT_RAM_05 = 256'hD0C937C9B730B4EA0520A1ED7A0400013C002130A7EAA1ED770400013C002151;
defparam dpb_inst_0.INIT_RAM_06 = 256'hFFBF309E30F433620040309EC930D431D90839000021EB08D9C9370228BB403E;
defparam dpb_inst_0.INIT_RAM_07 = 256'hC9F9C0BBFF3EE1C937D1335630F433625555309E30F43362AAAA309E30F43362;
defparam dpb_inst_0.INIT_RAM_08 = 256'h000801E1C90766FD066EFDC90566FD046EFDC9F9C0BB003EE1C9F9C0BB403EE1;
defparam dpb_inst_0.INIT_RAM_09 = 256'hD90839000021EB08D9C9F909FD000021FD0346FD024EFDC00186FD007EFD09FD;
defparam dpb_inst_0.INIT_RAM_0A = 256'h316131D90839000021EB08D93356FFF7347932C934443445310E345AC9314431;
defparam dpb_inst_0.INIT_RAM_0B = 256'h21031834F021053003CB08162F28BB2F2328BBFF3E316B200031B6347E3115C9;
defparam dpb_inst_0.INIT_RAM_0C = 256'hA1800031B634FA347DC93197311E18E52015318E200031B6347EC931863134EA;
defparam dpb_inst_0.INIT_RAM_0D = 256'h06373EC9FB20B1780BC1C9D9EBF9D931B1800031B634F6347DC931A7310E1831;
defparam dpb_inst_0.INIT_RAM_0E = 256'h08D9003E6F7DDD677CDDC9C1C9EE103D23DD2E0036DD04180077DD053003CB08;
defparam dpb_inst_0.INIT_RAM_0F = 256'hDD33563208010031D43E80345732B934443E583457C931EB31D90839000021EB;
defparam dpb_inst_0.INIT_RAM_10 = 256'h304333204D415256204B3120C93208EAA1ED23DD3C0077DD003E0400013C0021;
defparam dpb_inst_0.INIT_RAM_11 = 256'h204B36310020464646342D30303034204D415244204B34200020464646332D30;
defparam dpb_inst_0.INIT_RAM_12 = 256'h46422D30303038204D415244204B36310020464646372D30303034204D415244;
defparam dpb_inst_0.INIT_RAM_13 = 256'h4D2030382D5352540020464646462D30303043204D415244204B363100204646;
defparam dpb_inst_0.INIT_RAM_14 = 256'h202F20465744385A49204B4E415246202D2D204D4F52205453455420334D2F31;
defparam dpb_inst_0.INIT_RAM_15 = 256'h4341524148432D004B43414C42204E4149524441202F205633494B2045564144;
defparam dpb_inst_0.INIT_RAM_16 = 256'h54494200202D2D2D4B4F2D2D2D00202E2E545345542E2E002D54455320524554;
defparam dpb_inst_0.INIT_RAM_17 = 256'h2820214B4F002931204C45444F4D205449422D372820214B4F00205352524520;
defparam dpb_inst_0.INIT_RAM_18 = 256'h143C000400002020455A4953204B4E414220474E495453455400295449422D38;
defparam dpb_inst_0.INIT_RAM_19 = 256'h64C000400035063250800040003500323C40004000350033077000100034C632;
defparam dpb_inst_0.INIT_RAM_1A = 256'hD8E1C9F9E1C9D9EBF9D9C9E1FD334700003500322840001000332B0000351032;
defparam dpb_inst_0.INIT_RAM_1B = 256'h772F010E440366FD026EFD575FAFC9F9D90839000021EB08D9E1C9F9D0E1C9F9;
defparam dpb_inst_0.INIT_RAM_1C = 256'hB0790B23720366FD026EFD0146FD004EFD4D18FF1E0418F62800FE0628BE022F;
defparam dpb_inst_0.INIT_RAM_1D = 256'h4EFDF020B0790B23772F7A5FB3AA0428BA7E0366FD026EFD0146FD004EFDF920;
defparam dpb_inst_0.INIT_RAM_1E = 256'hAF1861180418F020B0790B23727A5FB3AA0428BA2F7E0366FD026EFD0146FD00;
defparam dpb_inst_0.INIT_RAM_1F = 256'h4EFDF020B0790B2B772F7A5FB3AA0428BA7E2B090366FD026EFD0146FD004EFD;
defparam dpb_inst_0.INIT_RAM_20 = 256'hFD004EFDF020B0790B2B727A5FB3AA0428BA2F7E2B090366FD026EFD0146FD00;
defparam dpb_inst_0.INIT_RAM_21 = 256'h979F28551600FE7AF220B0790B2B7A5FB3AA0428BA7E2B090366FD026EFD0146;
defparam dpb_inst_0.INIT_RAM_22 = 256'h40C6C0E67DDDC9E1DDC93C0021DDC9F4182323DD0077DD0828B77EE1C937C8B3;
defparam dpb_inst_0.INIT_RAM_23 = 256'h794EE1C909DDC1C93C0021DD346DEAA1ED20360400013C0021C924DD02306FDD;
defparam dpb_inst_0.INIT_RAM_24 = 256'h18FFD34603EEFC100018FFD34603EEFC100018FFD346023E2628B77E233A28B7;
defparam dpb_inst_0.INIT_RAM_25 = 256'hD3003EC118237EF5200DFA100018001800060B18DE200DE1204FCB03EEFC1000;
defparam dpb_inst_0.INIT_RAM_26 = 256'h9004A004B003C0030000C060501090105010901050109010501000004060C9FF;
defparam dpb_inst_0.INIT_RAM_27 = 256'h00000080C044000030FF00000020C01000000020304000005040600570058004;
defparam dpb_inst_0.INIT_RAM_28 = 256'h0000000000606040001060400010604000000060604000106040000000606040;

endmodule //Gowin_DPB2
