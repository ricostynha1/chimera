// This program was cloned from: https://github.com/neogeodev/NeoGeoFPGA-sim
// License: GNU General Public License v3.0

module jedi_lut (
	output reg [15:0] dout,
	input [13:0] address
);

	// Todo: dout could be only 12 bits ?

	always @(address)
	begin
		case (address)
		14'd0 : dout <=  16'd2;
		14'd1 : dout <=  16'd6;
		14'd2 : dout <=  16'd10;
		14'd3 : dout <=  16'd14;
		14'd4 : dout <=  16'd18;
		14'd5 : dout <=  16'd22;
		14'd6 : dout <=  16'd26;
		14'd7 : dout <=  16'd30;
		14'd8 : dout <= -16'd2;
		14'd9 : dout <= -16'd6;
		14'd10 : dout <= -16'd10;
		14'd11 : dout <= -16'd14;
		14'd12 : dout <= -16'd18;
		14'd13 : dout <= -16'd22;
		14'd14 : dout <= -16'd26;
		14'd15 : dout <= -16'd30;
		14'd16 : dout <=  16'd2;
		14'd17 : dout <=  16'd6;
		14'd18 : dout <=  16'd10;
		14'd19 : dout <=  16'd14;
		14'd20 : dout <=  16'd19;
		14'd21 : dout <=  16'd23;
		14'd22 : dout <=  16'd27;
		14'd23 : dout <=  16'd31;
		14'd24 : dout <= -16'd2;
		14'd25 : dout <= -16'd6;
		14'd26 : dout <= -16'd10;
		14'd27 : dout <= -16'd14;
		14'd28 : dout <= -16'd19;
		14'd29 : dout <= -16'd23;
		14'd30 : dout <= -16'd27;
		14'd31 : dout <= -16'd31;
		14'd32 : dout <=  16'd2;
		14'd33 : dout <=  16'd7;
		14'd34 : dout <=  16'd11;
		14'd35 : dout <=  16'd16;
		14'd36 : dout <=  16'd21;
		14'd37 : dout <=  16'd26;
		14'd38 : dout <=  16'd30;
		14'd39 : dout <=  16'd35;
		14'd40 : dout <= -16'd2;
		14'd41 : dout <= -16'd7;
		14'd42 : dout <= -16'd11;
		14'd43 : dout <= -16'd16;
		14'd44 : dout <= -16'd21;
		14'd45 : dout <= -16'd26;
		14'd46 : dout <= -16'd30;
		14'd47 : dout <= -16'd35;
		14'd48 : dout <=  16'd2;
		14'd49 : dout <=  16'd7;
		14'd50 : dout <=  16'd13;
		14'd51 : dout <=  16'd18;
		14'd52 : dout <=  16'd23;
		14'd53 : dout <=  16'd28;
		14'd54 : dout <=  16'd34;
		14'd55 : dout <=  16'd39;
		14'd56 : dout <= -16'd2;
		14'd57 : dout <= -16'd7;
		14'd58 : dout <= -16'd13;
		14'd59 : dout <= -16'd18;
		14'd60 : dout <= -16'd23;
		14'd61 : dout <= -16'd28;
		14'd62 : dout <= -16'd34;
		14'd63 : dout <= -16'd39;
		14'd64 : dout <=  16'd2;
		14'd65 : dout <=  16'd8;
		14'd66 : dout <=  16'd14;
		14'd67 : dout <=  16'd20;
		14'd68 : dout <=  16'd25;
		14'd69 : dout <=  16'd31;
		14'd70 : dout <=  16'd37;
		14'd71 : dout <=  16'd43;
		14'd72 : dout <= -16'd2;
		14'd73 : dout <= -16'd8;
		14'd74 : dout <= -16'd14;
		14'd75 : dout <= -16'd20;
		14'd76 : dout <= -16'd25;
		14'd77 : dout <= -16'd31;
		14'd78 : dout <= -16'd37;
		14'd79 : dout <= -16'd43;
		14'd80 : dout <=  16'd3;
		14'd81 : dout <=  16'd9;
		14'd82 : dout <=  16'd15;
		14'd83 : dout <=  16'd21;
		14'd84 : dout <=  16'd28;
		14'd85 : dout <=  16'd34;
		14'd86 : dout <=  16'd40;
		14'd87 : dout <=  16'd46;
		14'd88 : dout <= -16'd3;
		14'd89 : dout <= -16'd9;
		14'd90 : dout <= -16'd15;
		14'd91 : dout <= -16'd21;
		14'd92 : dout <= -16'd28;
		14'd93 : dout <= -16'd34;
		14'd94 : dout <= -16'd40;
		14'd95 : dout <= -16'd46;
		14'd96 : dout <=  16'd3;
		14'd97 : dout <=  16'd10;
		14'd98 : dout <=  16'd17;
		14'd99 : dout <=  16'd24;
		14'd100 : dout <=  16'd31;
		14'd101 : dout <=  16'd38;
		14'd102 : dout <=  16'd45;
		14'd103 : dout <=  16'd52;
		14'd104 : dout <= -16'd3;
		14'd105 : dout <= -16'd10;
		14'd106 : dout <= -16'd17;
		14'd107 : dout <= -16'd24;
		14'd108 : dout <= -16'd31;
		14'd109 : dout <= -16'd38;
		14'd110 : dout <= -16'd45;
		14'd111 : dout <= -16'd52;
		14'd112 : dout <=  16'd3;
		14'd113 : dout <=  16'd11;
		14'd114 : dout <=  16'd19;
		14'd115 : dout <=  16'd27;
		14'd116 : dout <=  16'd34;
		14'd117 : dout <=  16'd42;
		14'd118 : dout <=  16'd50;
		14'd119 : dout <=  16'd58;
		14'd120 : dout <= -16'd3;
		14'd121 : dout <= -16'd11;
		14'd122 : dout <= -16'd19;
		14'd123 : dout <= -16'd27;
		14'd124 : dout <= -16'd34;
		14'd125 : dout <= -16'd42;
		14'd126 : dout <= -16'd50;
		14'd127 : dout <= -16'd58;
		14'd128 : dout <=  16'd4;
		14'd129 : dout <=  16'd12;
		14'd130 : dout <=  16'd21;
		14'd131 : dout <=  16'd29;
		14'd132 : dout <=  16'd38;
		14'd133 : dout <=  16'd46;
		14'd134 : dout <=  16'd55;
		14'd135 : dout <=  16'd63;
		14'd136 : dout <= -16'd4;
		14'd137 : dout <= -16'd12;
		14'd138 : dout <= -16'd21;
		14'd139 : dout <= -16'd29;
		14'd140 : dout <= -16'd38;
		14'd141 : dout <= -16'd46;
		14'd142 : dout <= -16'd55;
		14'd143 : dout <= -16'd63;
		14'd144 : dout <=  16'd4;
		14'd145 : dout <=  16'd13;
		14'd146 : dout <=  16'd23;
		14'd147 : dout <=  16'd32;
		14'd148 : dout <=  16'd41;
		14'd149 : dout <=  16'd50;
		14'd150 : dout <=  16'd60;
		14'd151 : dout <=  16'd69;
		14'd152 : dout <= -16'd4;
		14'd153 : dout <= -16'd13;
		14'd154 : dout <= -16'd23;
		14'd155 : dout <= -16'd32;
		14'd156 : dout <= -16'd41;
		14'd157 : dout <= -16'd50;
		14'd158 : dout <= -16'd60;
		14'd159 : dout <= -16'd69;
		14'd160 : dout <=  16'd5;
		14'd161 : dout <=  16'd15;
		14'd162 : dout <=  16'd25;
		14'd163 : dout <=  16'd35;
		14'd164 : dout <=  16'd46;
		14'd165 : dout <=  16'd56;
		14'd166 : dout <=  16'd66;
		14'd167 : dout <=  16'd76;
		14'd168 : dout <= -16'd5;
		14'd169 : dout <= -16'd15;
		14'd170 : dout <= -16'd25;
		14'd171 : dout <= -16'd35;
		14'd172 : dout <= -16'd46;
		14'd173 : dout <= -16'd56;
		14'd174 : dout <= -16'd66;
		14'd175 : dout <= -16'd76;
		14'd176 : dout <=  16'd5;
		14'd177 : dout <=  16'd16;
		14'd178 : dout <=  16'd28;
		14'd179 : dout <=  16'd39;
		14'd180 : dout <=  16'd50;
		14'd181 : dout <=  16'd61;
		14'd182 : dout <=  16'd73;
		14'd183 : dout <=  16'd84;
		14'd184 : dout <= -16'd5;
		14'd185 : dout <= -16'd16;
		14'd186 : dout <= -16'd28;
		14'd187 : dout <= -16'd39;
		14'd188 : dout <= -16'd50;
		14'd189 : dout <= -16'd61;
		14'd190 : dout <= -16'd73;
		14'd191 : dout <= -16'd84;
		14'd192 : dout <=  16'd6;
		14'd193 : dout <=  16'd18;
		14'd194 : dout <=  16'd31;
		14'd195 : dout <=  16'd43;
		14'd196 : dout <=  16'd56;
		14'd197 : dout <=  16'd68;
		14'd198 : dout <=  16'd81;
		14'd199 : dout <=  16'd93;
		14'd200 : dout <= -16'd6;
		14'd201 : dout <= -16'd18;
		14'd202 : dout <= -16'd31;
		14'd203 : dout <= -16'd43;
		14'd204 : dout <= -16'd56;
		14'd205 : dout <= -16'd68;
		14'd206 : dout <= -16'd81;
		14'd207 : dout <= -16'd93;
		14'd208 : dout <=  16'd6;
		14'd209 : dout <=  16'd20;
		14'd210 : dout <=  16'd34;
		14'd211 : dout <=  16'd48;
		14'd212 : dout <=  16'd61;
		14'd213 : dout <=  16'd75;
		14'd214 : dout <=  16'd89;
		14'd215 : dout <=  16'd103;
		14'd216 : dout <= -16'd6;
		14'd217 : dout <= -16'd20;
		14'd218 : dout <= -16'd34;
		14'd219 : dout <= -16'd48;
		14'd220 : dout <= -16'd61;
		14'd221 : dout <= -16'd75;
		14'd222 : dout <= -16'd89;
		14'd223 : dout <= -16'd103;
		14'd224 : dout <=  16'd7;
		14'd225 : dout <=  16'd22;
		14'd226 : dout <=  16'd37;
		14'd227 : dout <=  16'd52;
		14'd228 : dout <=  16'd67;
		14'd229 : dout <=  16'd82;
		14'd230 : dout <=  16'd97;
		14'd231 : dout <=  16'd112;
		14'd232 : dout <= -16'd7;
		14'd233 : dout <= -16'd22;
		14'd234 : dout <= -16'd37;
		14'd235 : dout <= -16'd52;
		14'd236 : dout <= -16'd67;
		14'd237 : dout <= -16'd82;
		14'd238 : dout <= -16'd97;
		14'd239 : dout <= -16'd112;
		14'd240 : dout <=  16'd8;
		14'd241 : dout <=  16'd24;
		14'd242 : dout <=  16'd41;
		14'd243 : dout <=  16'd57;
		14'd244 : dout <=  16'd74;
		14'd245 : dout <=  16'd90;
		14'd246 : dout <=  16'd107;
		14'd247 : dout <=  16'd123;
		14'd248 : dout <= -16'd8;
		14'd249 : dout <= -16'd24;
		14'd250 : dout <= -16'd41;
		14'd251 : dout <= -16'd57;
		14'd252 : dout <= -16'd74;
		14'd253 : dout <= -16'd90;
		14'd254 : dout <= -16'd107;
		14'd255 : dout <= -16'd123;
		14'd256 : dout <=  16'd9;
		14'd257 : dout <=  16'd27;
		14'd258 : dout <=  16'd45;
		14'd259 : dout <=  16'd63;
		14'd260 : dout <=  16'd82;
		14'd261 : dout <=  16'd100;
		14'd262 : dout <=  16'd118;
		14'd263 : dout <=  16'd136;
		14'd264 : dout <= -16'd9;
		14'd265 : dout <= -16'd27;
		14'd266 : dout <= -16'd45;
		14'd267 : dout <= -16'd63;
		14'd268 : dout <= -16'd82;
		14'd269 : dout <= -16'd100;
		14'd270 : dout <= -16'd118;
		14'd271 : dout <= -16'd136;
		14'd272 : dout <=  16'd10;
		14'd273 : dout <=  16'd30;
		14'd274 : dout <=  16'd50;
		14'd275 : dout <=  16'd70;
		14'd276 : dout <=  16'd90;
		14'd277 : dout <=  16'd110;
		14'd278 : dout <=  16'd130;
		14'd279 : dout <=  16'd150;
		14'd280 : dout <= -16'd10;
		14'd281 : dout <= -16'd30;
		14'd282 : dout <= -16'd50;
		14'd283 : dout <= -16'd70;
		14'd284 : dout <= -16'd90;
		14'd285 : dout <= -16'd110;
		14'd286 : dout <= -16'd130;
		14'd287 : dout <= -16'd150;
		14'd288 : dout <=  16'd11;
		14'd289 : dout <=  16'd33;
		14'd290 : dout <=  16'd55;
		14'd291 : dout <=  16'd77;
		14'd292 : dout <=  16'd99;
		14'd293 : dout <=  16'd121;
		14'd294 : dout <=  16'd143;
		14'd295 : dout <=  16'd165;
		14'd296 : dout <= -16'd11;
		14'd297 : dout <= -16'd33;
		14'd298 : dout <= -16'd55;
		14'd299 : dout <= -16'd77;
		14'd300 : dout <= -16'd99;
		14'd301 : dout <= -16'd121;
		14'd302 : dout <= -16'd143;
		14'd303 : dout <= -16'd165;
		14'd304 : dout <=  16'd12;
		14'd305 : dout <=  16'd36;
		14'd306 : dout <=  16'd60;
		14'd307 : dout <=  16'd84;
		14'd308 : dout <=  16'd109;
		14'd309 : dout <=  16'd133;
		14'd310 : dout <=  16'd157;
		14'd311 : dout <=  16'd181;
		14'd312 : dout <= -16'd12;
		14'd313 : dout <= -16'd36;
		14'd314 : dout <= -16'd60;
		14'd315 : dout <= -16'd84;
		14'd316 : dout <= -16'd109;
		14'd317 : dout <= -16'd133;
		14'd318 : dout <= -16'd157;
		14'd319 : dout <= -16'd181;
		14'd320 : dout <=  16'd13;
		14'd321 : dout <=  16'd40;
		14'd322 : dout <=  16'd66;
		14'd323 : dout <=  16'd93;
		14'd324 : dout <=  16'd120;
		14'd325 : dout <=  16'd147;
		14'd326 : dout <=  16'd173;
		14'd327 : dout <=  16'd200;
		14'd328 : dout <= -16'd13;
		14'd329 : dout <= -16'd40;
		14'd330 : dout <= -16'd66;
		14'd331 : dout <= -16'd93;
		14'd332 : dout <= -16'd120;
		14'd333 : dout <= -16'd147;
		14'd334 : dout <= -16'd173;
		14'd335 : dout <= -16'd200;
		14'd336 : dout <=  16'd14;
		14'd337 : dout <=  16'd44;
		14'd338 : dout <=  16'd73;
		14'd339 : dout <=  16'd103;
		14'd340 : dout <=  16'd132;
		14'd341 : dout <=  16'd162;
		14'd342 : dout <=  16'd191;
		14'd343 : dout <=  16'd221;
		14'd344 : dout <= -16'd14;
		14'd345 : dout <= -16'd44;
		14'd346 : dout <= -16'd73;
		14'd347 : dout <= -16'd103;
		14'd348 : dout <= -16'd132;
		14'd349 : dout <= -16'd162;
		14'd350 : dout <= -16'd191;
		14'd351 : dout <= -16'd221;
		14'd352 : dout <=  16'd16;
		14'd353 : dout <=  16'd48;
		14'd354 : dout <=  16'd81;
		14'd355 : dout <=  16'd113;
		14'd356 : dout <=  16'd146;
		14'd357 : dout <=  16'd178;
		14'd358 : dout <=  16'd211;
		14'd359 : dout <=  16'd243;
		14'd360 : dout <= -16'd16;
		14'd361 : dout <= -16'd48;
		14'd362 : dout <= -16'd81;
		14'd363 : dout <= -16'd113;
		14'd364 : dout <= -16'd146;
		14'd365 : dout <= -16'd178;
		14'd366 : dout <= -16'd211;
		14'd367 : dout <= -16'd243;
		14'd368 : dout <=  16'd17;
		14'd369 : dout <=  16'd53;
		14'd370 : dout <=  16'd89;
		14'd371 : dout <=  16'd125;
		14'd372 : dout <=  16'd160;
		14'd373 : dout <=  16'd196;
		14'd374 : dout <=  16'd232;
		14'd375 : dout <=  16'd268;
		14'd376 : dout <= -16'd17;
		14'd377 : dout <= -16'd53;
		14'd378 : dout <= -16'd89;
		14'd379 : dout <= -16'd125;
		14'd380 : dout <= -16'd160;
		14'd381 : dout <= -16'd196;
		14'd382 : dout <= -16'd232;
		14'd383 : dout <= -16'd268;
		14'd384 : dout <=  16'd19;
		14'd385 : dout <=  16'd58;
		14'd386 : dout <=  16'd98;
		14'd387 : dout <=  16'd137;
		14'd388 : dout <=  16'd176;
		14'd389 : dout <=  16'd215;
		14'd390 : dout <=  16'd255;
		14'd391 : dout <=  16'd294;
		14'd392 : dout <= -16'd19;
		14'd393 : dout <= -16'd58;
		14'd394 : dout <= -16'd98;
		14'd395 : dout <= -16'd137;
		14'd396 : dout <= -16'd176;
		14'd397 : dout <= -16'd215;
		14'd398 : dout <= -16'd255;
		14'd399 : dout <= -16'd294;
		14'd400 : dout <=  16'd21;
		14'd401 : dout <=  16'd64;
		14'd402 : dout <=  16'd108;
		14'd403 : dout <=  16'd151;
		14'd404 : dout <=  16'd194;
		14'd405 : dout <=  16'd237;
		14'd406 : dout <=  16'd281;
		14'd407 : dout <=  16'd324;
		14'd408 : dout <= -16'd21;
		14'd409 : dout <= -16'd64;
		14'd410 : dout <= -16'd108;
		14'd411 : dout <= -16'd151;
		14'd412 : dout <= -16'd194;
		14'd413 : dout <= -16'd237;
		14'd414 : dout <= -16'd281;
		14'd415 : dout <= -16'd324;
		14'd416 : dout <=  16'd23;
		14'd417 : dout <=  16'd71;
		14'd418 : dout <=  16'd118;
		14'd419 : dout <=  16'd166;
		14'd420 : dout <=  16'd213;
		14'd421 : dout <=  16'd261;
		14'd422 : dout <=  16'd308;
		14'd423 : dout <=  16'd356;
		14'd424 : dout <= -16'd23;
		14'd425 : dout <= -16'd71;
		14'd426 : dout <= -16'd118;
		14'd427 : dout <= -16'd166;
		14'd428 : dout <= -16'd213;
		14'd429 : dout <= -16'd261;
		14'd430 : dout <= -16'd308;
		14'd431 : dout <= -16'd356;
		14'd432 : dout <=  16'd26;
		14'd433 : dout <=  16'd78;
		14'd434 : dout <=  16'd130;
		14'd435 : dout <=  16'd182;
		14'd436 : dout <=  16'd235;
		14'd437 : dout <=  16'd287;
		14'd438 : dout <=  16'd339;
		14'd439 : dout <=  16'd391;
		14'd440 : dout <= -16'd26;
		14'd441 : dout <= -16'd78;
		14'd442 : dout <= -16'd130;
		14'd443 : dout <= -16'd182;
		14'd444 : dout <= -16'd235;
		14'd445 : dout <= -16'd287;
		14'd446 : dout <= -16'd339;
		14'd447 : dout <= -16'd391;
		14'd448 : dout <=  16'd28;
		14'd449 : dout <=  16'd86;
		14'd450 : dout <=  16'd143;
		14'd451 : dout <=  16'd201;
		14'd452 : dout <=  16'd258;
		14'd453 : dout <=  16'd316;
		14'd454 : dout <=  16'd373;
		14'd455 : dout <=  16'd431;
		14'd456 : dout <= -16'd28;
		14'd457 : dout <= -16'd86;
		14'd458 : dout <= -16'd143;
		14'd459 : dout <= -16'd201;
		14'd460 : dout <= -16'd258;
		14'd461 : dout <= -16'd316;
		14'd462 : dout <= -16'd373;
		14'd463 : dout <= -16'd431;
		14'd464 : dout <=  16'd31;
		14'd465 : dout <=  16'd94;
		14'd466 : dout <=  16'd158;
		14'd467 : dout <=  16'd221;
		14'd468 : dout <=  16'd284;
		14'd469 : dout <=  16'd347;
		14'd470 : dout <=  16'd411;
		14'd471 : dout <=  16'd474;
		14'd472 : dout <= -16'd31;
		14'd473 : dout <= -16'd94;
		14'd474 : dout <= -16'd158;
		14'd475 : dout <= -16'd221;
		14'd476 : dout <= -16'd284;
		14'd477 : dout <= -16'd347;
		14'd478 : dout <= -16'd411;
		14'd479 : dout <= -16'd474;
		14'd480 : dout <=  16'd34;
		14'd481 : dout <=  16'd104;
		14'd482 : dout <=  16'd174;
		14'd483 : dout <=  16'd244;
		14'd484 : dout <=  16'd313;
		14'd485 : dout <=  16'd383;
		14'd486 : dout <=  16'd453;
		14'd487 : dout <=  16'd523;
		14'd488 : dout <= -16'd34;
		14'd489 : dout <= -16'd104;
		14'd490 : dout <= -16'd174;
		14'd491 : dout <= -16'd244;
		14'd492 : dout <= -16'd313;
		14'd493 : dout <= -16'd383;
		14'd494 : dout <= -16'd453;
		14'd495 : dout <= -16'd523;
		14'd496 : dout <=  16'd38;
		14'd497 : dout <=  16'd115;
		14'd498 : dout <=  16'd191;
		14'd499 : dout <=  16'd268;
		14'd500 : dout <=  16'd345;
		14'd501 : dout <=  16'd422;
		14'd502 : dout <=  16'd498;
		14'd503 : dout <=  16'd575;
		14'd504 : dout <= -16'd38;
		14'd505 : dout <= -16'd115;
		14'd506 : dout <= -16'd191;
		14'd507 : dout <= -16'd268;
		14'd508 : dout <= -16'd345;
		14'd509 : dout <= -16'd422;
		14'd510 : dout <= -16'd498;
		14'd511 : dout <= -16'd575;
		14'd512 : dout <=  16'd42;
		14'd513 : dout <=  16'd126;
		14'd514 : dout <=  16'd210;
		14'd515 : dout <=  16'd294;
		14'd516 : dout <=  16'd379;
		14'd517 : dout <=  16'd463;
		14'd518 : dout <=  16'd547;
		14'd519 : dout <=  16'd631;
		14'd520 : dout <= -16'd42;
		14'd521 : dout <= -16'd126;
		14'd522 : dout <= -16'd210;
		14'd523 : dout <= -16'd294;
		14'd524 : dout <= -16'd379;
		14'd525 : dout <= -16'd463;
		14'd526 : dout <= -16'd547;
		14'd527 : dout <= -16'd631;
		14'd528 : dout <=  16'd46;
		14'd529 : dout <=  16'd139;
		14'd530 : dout <=  16'd231;
		14'd531 : dout <=  16'd324;
		14'd532 : dout <=  16'd417;
		14'd533 : dout <=  16'd510;
		14'd534 : dout <=  16'd602;
		14'd535 : dout <=  16'd695;
		14'd536 : dout <= -16'd46;
		14'd537 : dout <= -16'd139;
		14'd538 : dout <= -16'd231;
		14'd539 : dout <= -16'd324;
		14'd540 : dout <= -16'd417;
		14'd541 : dout <= -16'd510;
		14'd542 : dout <= -16'd602;
		14'd543 : dout <= -16'd695;
		14'd544 : dout <=  16'd51;
		14'd545 : dout <=  16'd153;
		14'd546 : dout <=  16'd255;
		14'd547 : dout <=  16'd357;
		14'd548 : dout <=  16'd459;
		14'd549 : dout <=  16'd561;
		14'd550 : dout <=  16'd663;
		14'd551 : dout <=  16'd765;
		14'd552 : dout <= -16'd51;
		14'd553 : dout <= -16'd153;
		14'd554 : dout <= -16'd255;
		14'd555 : dout <= -16'd357;
		14'd556 : dout <= -16'd459;
		14'd557 : dout <= -16'd561;
		14'd558 : dout <= -16'd663;
		14'd559 : dout <= -16'd765;
		14'd560 : dout <=  16'd56;
		14'd561 : dout <=  16'd168;
		14'd562 : dout <=  16'd280;
		14'd563 : dout <=  16'd392;
		14'd564 : dout <=  16'd505;
		14'd565 : dout <=  16'd617;
		14'd566 : dout <=  16'd729;
		14'd567 : dout <=  16'd841;
		14'd568 : dout <= -16'd56;
		14'd569 : dout <= -16'd168;
		14'd570 : dout <= -16'd280;
		14'd571 : dout <= -16'd392;
		14'd572 : dout <= -16'd505;
		14'd573 : dout <= -16'd617;
		14'd574 : dout <= -16'd729;
		14'd575 : dout <= -16'd841;
		14'd576 : dout <=  16'd61;
		14'd577 : dout <=  16'd185;
		14'd578 : dout <=  16'd308;
		14'd579 : dout <=  16'd432;
		14'd580 : dout <=  16'd555;
		14'd581 : dout <=  16'd679;
		14'd582 : dout <=  16'd802;
		14'd583 : dout <=  16'd926;
		14'd584 : dout <= -16'd61;
		14'd585 : dout <= -16'd185;
		14'd586 : dout <= -16'd308;
		14'd587 : dout <= -16'd432;
		14'd588 : dout <= -16'd555;
		14'd589 : dout <= -16'd679;
		14'd590 : dout <= -16'd802;
		14'd591 : dout <= -16'd926;
		14'd592 : dout <=  16'd68;
		14'd593 : dout <=  16'd204;
		14'd594 : dout <=  16'd340;
		14'd595 : dout <=  16'd476;
		14'd596 : dout <=  16'd612;
		14'd597 : dout <=  16'd748;
		14'd598 : dout <=  16'd884;
		14'd599 : dout <=  16'd1020;
		14'd600 : dout <= -16'd68;
		14'd601 : dout <= -16'd204;
		14'd602 : dout <= -16'd340;
		14'd603 : dout <= -16'd476;
		14'd604 : dout <= -16'd612;
		14'd605 : dout <= -16'd748;
		14'd606 : dout <= -16'd884;
		14'd607 : dout <= -16'd1020;
		14'd608 : dout <=  16'd74;
		14'd609 : dout <=  16'd224;
		14'd610 : dout <=  16'd373;
		14'd611 : dout <=  16'd523;
		14'd612 : dout <=  16'd672;
		14'd613 : dout <=  16'd822;
		14'd614 : dout <=  16'd971;
		14'd615 : dout <=  16'd1121;
		14'd616 : dout <= -16'd74;
		14'd617 : dout <= -16'd224;
		14'd618 : dout <= -16'd373;
		14'd619 : dout <= -16'd523;
		14'd620 : dout <= -16'd672;
		14'd621 : dout <= -16'd822;
		14'd622 : dout <= -16'd971;
		14'd623 : dout <= -16'd1121;
		14'd624 : dout <=  16'd82;
		14'd625 : dout <=  16'd246;
		14'd626 : dout <=  16'd411;
		14'd627 : dout <=  16'd575;
		14'd628 : dout <=  16'd740;
		14'd629 : dout <=  16'd904;
		14'd630 : dout <=  16'd1069;
		14'd631 : dout <=  16'd1233;
		14'd632 : dout <= -16'd82;
		14'd633 : dout <= -16'd246;
		14'd634 : dout <= -16'd411;
		14'd635 : dout <= -16'd575;
		14'd636 : dout <= -16'd740;
		14'd637 : dout <= -16'd904;
		14'd638 : dout <= -16'd1069;
		14'd639 : dout <= -16'd1233;
		14'd640 : dout <=  16'd90;
		14'd641 : dout <=  16'd271;
		14'd642 : dout <=  16'd452;
		14'd643 : dout <=  16'd633;
		14'd644 : dout <=  16'd814;
		14'd645 : dout <=  16'd995;
		14'd646 : dout <=  16'd1176;
		14'd647 : dout <=  16'd1357;
		14'd648 : dout <= -16'd90;
		14'd649 : dout <= -16'd271;
		14'd650 : dout <= -16'd452;
		14'd651 : dout <= -16'd633;
		14'd652 : dout <= -16'd814;
		14'd653 : dout <= -16'd995;
		14'd654 : dout <= -16'd1176;
		14'd655 : dout <= -16'd1357;
		14'd656 : dout <=  16'd99;
		14'd657 : dout <=  16'd298;
		14'd658 : dout <=  16'd497;
		14'd659 : dout <=  16'd696;
		14'd660 : dout <=  16'd895;
		14'd661 : dout <=  16'd1094;
		14'd662 : dout <=  16'd1293;
		14'd663 : dout <=  16'd1492;
		14'd664 : dout <= -16'd99;
		14'd665 : dout <= -16'd298;
		14'd666 : dout <= -16'd497;
		14'd667 : dout <= -16'd696;
		14'd668 : dout <= -16'd895;
		14'd669 : dout <= -16'd1094;
		14'd670 : dout <= -16'd1293;
		14'd671 : dout <= -16'd1492;
		14'd672 : dout <=  16'd109;
		14'd673 : dout <=  16'd328;
		14'd674 : dout <=  16'd547;
		14'd675 : dout <=  16'd766;
		14'd676 : dout <=  16'd985;
		14'd677 : dout <=  16'd1204;
		14'd678 : dout <=  16'd1423;
		14'd679 : dout <=  16'd1642;
		14'd680 : dout <= -16'd109;
		14'd681 : dout <= -16'd328;
		14'd682 : dout <= -16'd547;
		14'd683 : dout <= -16'd766;
		14'd684 : dout <= -16'd985;
		14'd685 : dout <= -16'd1204;
		14'd686 : dout <= -16'd1423;
		14'd687 : dout <= -16'd1642;
		14'd688 : dout <=  16'd120;
		14'd689 : dout <=  16'd361;
		14'd690 : dout <=  16'd601;
		14'd691 : dout <=  16'd842;
		14'd692 : dout <=  16'd1083;
		14'd693 : dout <=  16'd1324;
		14'd694 : dout <=  16'd1564;
		14'd695 : dout <=  16'd1805;
		14'd696 : dout <= -16'd120;
		14'd697 : dout <= -16'd361;
		14'd698 : dout <= -16'd601;
		14'd699 : dout <= -16'd842;
		14'd700 : dout <= -16'd1083;
		14'd701 : dout <= -16'd1324;
		14'd702 : dout <= -16'd1564;
		14'd703 : dout <= -16'd1805;
		14'd704 : dout <=  16'd132;
		14'd705 : dout <=  16'd397;
		14'd706 : dout <=  16'd662;
		14'd707 : dout <=  16'd927;
		14'd708 : dout <=  16'd1192;
		14'd709 : dout <=  16'd1457;
		14'd710 : dout <=  16'd1722;
		14'd711 : dout <=  16'd1987;
		14'd712 : dout <= -16'd132;
		14'd713 : dout <= -16'd397;
		14'd714 : dout <= -16'd662;
		14'd715 : dout <= -16'd927;
		14'd716 : dout <= -16'd1192;
		14'd717 : dout <= -16'd1457;
		14'd718 : dout <= -16'd1722;
		14'd719 : dout <= -16'd1987;
		14'd720 : dout <=  16'd145;
		14'd721 : dout <=  16'd437;
		14'd722 : dout <=  16'd728;
		14'd723 : dout <=  16'd1020;
		14'd724 : dout <=  16'd1311;
		14'd725 : dout <=  16'd1603;
		14'd726 : dout <=  16'd1894;
		14'd727 : dout <=  16'd2186;
		14'd728 : dout <= -16'd145;
		14'd729 : dout <= -16'd437;
		14'd730 : dout <= -16'd728;
		14'd731 : dout <= -16'd1020;
		14'd732 : dout <= -16'd1311;
		14'd733 : dout <= -16'd1603;
		14'd734 : dout <= -16'd1894;
		14'd735 : dout <= -16'd2186;
		14'd736 : dout <=  16'd160;
		14'd737 : dout <=  16'd480;
		14'd738 : dout <=  16'd801;
		14'd739 : dout <=  16'd1121;
		14'd740 : dout <=  16'd1442;
		14'd741 : dout <=  16'd1762;
		14'd742 : dout <=  16'd2083;
		14'd743 : dout <=  16'd2403;
		14'd744 : dout <= -16'd160;
		14'd745 : dout <= -16'd480;
		14'd746 : dout <= -16'd801;
		14'd747 : dout <= -16'd1121;
		14'd748 : dout <= -16'd1442;
		14'd749 : dout <= -16'd1762;
		14'd750 : dout <= -16'd2083;
		14'd751 : dout <= -16'd2403;
		14'd752 : dout <=  16'd176;
		14'd753 : dout <=  16'd529;
		14'd754 : dout <=  16'd881;
		14'd755 : dout <=  16'd1234;
		14'd756 : dout <=  16'd1587;
		14'd757 : dout <=  16'd1940;
		14'd758 : dout <=  16'd2292;
		14'd759 : dout <=  16'd2645;
		14'd760 : dout <= -16'd176;
		14'd761 : dout <= -16'd529;
		14'd762 : dout <= -16'd881;
		14'd763 : dout <= -16'd1234;
		14'd764 : dout <= -16'd1587;
		14'd765 : dout <= -16'd1940;
		14'd766 : dout <= -16'd2292;
		14'd767 : dout <= -16'd2645;
		14'd768 : dout <=  16'd194;
		14'd769 : dout <=  16'd582;
		14'd770 : dout <=  16'd970;
		14'd771 : dout <=  16'd1358;
		14'd772 : dout <=  16'd1746;
		14'd773 : dout <=  16'd2134;
		14'd774 : dout <=  16'd2522;
		14'd775 : dout <=  16'd2910;
		14'd776 : dout <= -16'd194;
		14'd777 : dout <= -16'd582;
		14'd778 : dout <= -16'd970;
		14'd779 : dout <= -16'd1358;
		14'd780 : dout <= -16'd1746;
		14'd781 : dout <= -16'd2134;
		14'd782 : dout <= -16'd2522;
		14'd783 : dout <= -16'd2910;
		default : dout <= 16'd0;
		endcase
	end

endmodule
