// This program was cloned from: https://github.com/FIUSCIS-CDA/CPU_MultiCycle
// License: MIT License

///////////////////////////////////////////////////////////////////////////////////
// Component: MicroROM
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// Extended By: CDA3102 students
// License: MIT, (C) 2020-2022 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////

module MicroROM(state, microinstruction);
///////////////////////////////////////////////////////////////////////////////////
// Input: state (4-bit)
  input [4:0] state; 
///////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////
// Output: microinstruction (18-bit)
  output wire [19:0] microinstruction;
///////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////
// Internal: ROM
  reg [19:0] ROM[16:0];
///////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////
  // PUT MICROINSTRUCTIONS HERE
  // Bit Order: PCWrite, PCWriteCond, IorD, MemWrite, IRWrite, MemToReg (2),
  //            PCSrc (2), ALUOp (3), ALUSrcB (2), ALUSrcA, RegWrite,
  //            RegDst, isBNE, LOWrite, Shift16
  //////////////////////////////////////////////////////////////////////
  initial begin
  ROM[5'b00000] = 		20'b10001000000001000000;	// State 0
  ROM[5'b00001] =		20'b00000000000011000000;	// State 1
  ROM[5'b00010] =		20'b00000000000010100000;	// State 2
  ROM[5'b00011] =		20'b00100000000000000000; 	// State 3
  ROM[5'b00100] =		20'b00000010000000010000;	// State 4
  ROM[5'b00101] =		20'b00110000000000000000;	// State 5
  ROM[5'b00110] =		20'b00000000001000100000; 	// State 6
  ROM[5'b00111] = 		20'b00000000000000011000; 	// State 7
  ROM[5'b01000] = 		20'b01000000100100100000;	// State 8
  ROM[5'b01001] = 		20'b10000001000000000000;	// State 9
  ROM[5'b01010] =	     	20'b00000000000000010000;	// State 10
  ROM[5'b01011] =               20'b01000000100100100100; 	// State 11
  ROM[5'b01100] =               20'b00000000001110100000; 	// State 12  
  ROM[5'b01101] =               20'b00000000000000000010; 	// State 13
  ROM[5'b01110] =               20'b00000100000000011000; 	// State 14
  ROM[5'b01111] =               20'b00000000010010000001; 	// State 15
  ROM[5'b10000] =               20'b00000000010110100000; 	// State 16
  ////////////////////////////////////////////////////////////////////////
  end

  ////////////////////////////////////////////////////////////////////////
  // Microinstruction stored in ROM, address is the state
  assign microinstruction = ROM[state];
  ////////////////////////////////////////////////////////////////////////

endmodule
