// This program was cloned from: https://github.com/Nilesh002/Multiplication-and-Accumulation-Unit-MAC-
// License: MIT License

module add12(a,b,s);
input [11:0]a,b;
output [11:0]s;

assign s=a+b;

endmodule
