// This program was cloned from: https://github.com/rupin-r/CollegeProjects
// License: MIT License

module Design(input clock, input inputSerial, input reset, input uart_clock1, input uart_clock2, output [31:0] dataOut, output clkOut, output latch, output latch2, output clkCompare, output clkCompare2);
	
	reg [7:0] phase [255:0];
	reg [18:0] cnt;
	wire [255:0] select;
	reg [7:0] phase_end [255:0];
	wire [255:0] select_end;
	wire [255:0] values;
	reg [2:0] counter;
	reg [6:0] phase_count;
	reg [7:0] phase_edit;
	wire phase_clock;
	wire uart_clock;
	wire [7:0] newPhase;
	
	initial begin
		cnt = 0;
		//initial phases held in a pwm file that can be generated from the python code
		$readmemh("C:/altera/13.0sp1/quartus/pwm.txt", phase);
		counter = 0;
		phase_count = 0;
		phase_edit = 0;
	end
	
	//clock divider held in count
	always @(posedge clock) begin
		cnt = cnt + 1;
	end
	
	//responsible for shifting bits out
	always @(posedge cnt[0]) begin
		counter = counter + 1;
	end

	//turns on or off the bit based on whether the phase matches
	always @(posedge cnt[3]) begin
		phase_count = (phase_count + 1);
		if(phase_count == 80) begin
			phase_count = 0;
		end
	end	
	
	//edits the phases using UART communication
	UART_Receiver u(.clk(uart_clock), .rst_n(reset), .rx(inputSerial), .data(newPhase), .clkout(clkCompare));
	
	//takes the clock from the uart module that goes high only when receiving a full 8-bit phase to edit a phase
	always @(posedge clkCompare) begin
		//edit phases in order, loops back around after 255 since phase_edit is 8-bits
		phase[phase_edit] = newPhase;
		//adjust phase_end based on the following logic
			//phase_end = (phase + 40) % 80;
		//mod took too many resources so the logic was broken down as below:
		if(newPhase >= 40) begin
			phase_end[phase_edit] = newPhase - 40;
		end
		else begin
			phase_end[phase_edit] = newPhase + 40;
		end
		//increment the phase to edit
		phase_edit = phase_edit + 1;
	end
	
	//a clock signal that is high for 40 main clock signals and low for 40 main clock signals
	assign phase_clock = (phase_count[5] & (phase_count[4] || phase_count[3])) || phase_count[6];
	
	
	//each line follows the structure below, only changing the value [0] 
	//assign select[0] = (phase_count[0] ^ phase[0][0]) || (phase_count[1] ^ phase[0][1]) || (phase_count[2] ^ phase[0][2]) || (phase_count[3] ^ phase[0][3]) || (phase_count[4] ^ phase[0][4]) || (phase_count[5] ^ phase[0][5]) || (phase_count[6] ^ phase[0][6]) || phase[0][7];
	//logic is: select = 1 if MSB of phase is 1 or if select does not equal the phase of its emitter
	
	assign select[0] = (phase_count[0] ^ phase[0][0]) || (phase_count[1] ^ phase[0][1]) || (phase_count[2] ^ phase[0][2]) || (phase_count[3] ^ phase[0][3]) || (phase_count[4] ^ phase[0][4]) || (phase_count[5] ^ phase[0][5]) || (phase_count[6] ^ phase[0][6]) || phase[0][7];
	assign select[1] = (phase_count[0] ^ phase[1][0]) || (phase_count[1] ^ phase[1][1]) || (phase_count[2] ^ phase[1][2]) || (phase_count[3] ^ phase[1][3]) || (phase_count[4] ^ phase[1][4]) || (phase_count[5] ^ phase[1][5]) || (phase_count[6] ^ phase[1][6]) || phase[1][7];
	assign select[2] = (phase_count[0] ^ phase[2][0]) || (phase_count[1] ^ phase[2][1]) || (phase_count[2] ^ phase[2][2]) || (phase_count[3] ^ phase[2][3]) || (phase_count[4] ^ phase[2][4]) || (phase_count[5] ^ phase[2][5]) || (phase_count[6] ^ phase[2][6]) || phase[2][7];
	assign select[3] = (phase_count[0] ^ phase[3][0]) || (phase_count[1] ^ phase[3][1]) || (phase_count[2] ^ phase[3][2]) || (phase_count[3] ^ phase[3][3]) || (phase_count[4] ^ phase[3][4]) || (phase_count[5] ^ phase[3][5]) || (phase_count[6] ^ phase[3][6]) || phase[3][7];
	assign select[4] = (phase_count[0] ^ phase[4][0]) || (phase_count[1] ^ phase[4][1]) || (phase_count[2] ^ phase[4][2]) || (phase_count[3] ^ phase[4][3]) || (phase_count[4] ^ phase[4][4]) || (phase_count[5] ^ phase[4][5]) || (phase_count[6] ^ phase[4][6]) || phase[4][7];
	assign select[5] = (phase_count[0] ^ phase[5][0]) || (phase_count[1] ^ phase[5][1]) || (phase_count[2] ^ phase[5][2]) || (phase_count[3] ^ phase[5][3]) || (phase_count[4] ^ phase[5][4]) || (phase_count[5] ^ phase[5][5]) || (phase_count[6] ^ phase[5][6]) || phase[5][7];
	assign select[6] = (phase_count[0] ^ phase[6][0]) || (phase_count[1] ^ phase[6][1]) || (phase_count[2] ^ phase[6][2]) || (phase_count[3] ^ phase[6][3]) || (phase_count[4] ^ phase[6][4]) || (phase_count[5] ^ phase[6][5]) || (phase_count[6] ^ phase[6][6]) || phase[6][7];
	assign select[7] = (phase_count[0] ^ phase[7][0]) || (phase_count[1] ^ phase[7][1]) || (phase_count[2] ^ phase[7][2]) || (phase_count[3] ^ phase[7][3]) || (phase_count[4] ^ phase[7][4]) || (phase_count[5] ^ phase[7][5]) || (phase_count[6] ^ phase[7][6]) || phase[7][7];
	assign select[8] = (phase_count[0] ^ phase[8][0]) || (phase_count[1] ^ phase[8][1]) || (phase_count[2] ^ phase[8][2]) || (phase_count[3] ^ phase[8][3]) || (phase_count[4] ^ phase[8][4]) || (phase_count[5] ^ phase[8][5]) || (phase_count[6] ^ phase[8][6]) || phase[8][7];
	assign select[9] = (phase_count[0] ^ phase[9][0]) || (phase_count[1] ^ phase[9][1]) || (phase_count[2] ^ phase[9][2]) || (phase_count[3] ^ phase[9][3]) || (phase_count[4] ^ phase[9][4]) || (phase_count[5] ^ phase[9][5]) || (phase_count[6] ^ phase[9][6]) || phase[9][7];
	assign select[10] = (phase_count[0] ^ phase[10][0]) || (phase_count[1] ^ phase[10][1]) || (phase_count[2] ^ phase[10][2]) || (phase_count[3] ^ phase[10][3]) || (phase_count[4] ^ phase[10][4]) || (phase_count[5] ^ phase[10][5]) || (phase_count[6] ^ phase[10][6]) || phase[10][7];
	assign select[11] = (phase_count[0] ^ phase[11][0]) || (phase_count[1] ^ phase[11][1]) || (phase_count[2] ^ phase[11][2]) || (phase_count[3] ^ phase[11][3]) || (phase_count[4] ^ phase[11][4]) || (phase_count[5] ^ phase[11][5]) || (phase_count[6] ^ phase[11][6]) || phase[11][7];
	assign select[12] = (phase_count[0] ^ phase[12][0]) || (phase_count[1] ^ phase[12][1]) || (phase_count[2] ^ phase[12][2]) || (phase_count[3] ^ phase[12][3]) || (phase_count[4] ^ phase[12][4]) || (phase_count[5] ^ phase[12][5]) || (phase_count[6] ^ phase[12][6]) || phase[12][7];
	assign select[13] = (phase_count[0] ^ phase[13][0]) || (phase_count[1] ^ phase[13][1]) || (phase_count[2] ^ phase[13][2]) || (phase_count[3] ^ phase[13][3]) || (phase_count[4] ^ phase[13][4]) || (phase_count[5] ^ phase[13][5]) || (phase_count[6] ^ phase[13][6]) || phase[13][7];
	assign select[14] = (phase_count[0] ^ phase[14][0]) || (phase_count[1] ^ phase[14][1]) || (phase_count[2] ^ phase[14][2]) || (phase_count[3] ^ phase[14][3]) || (phase_count[4] ^ phase[14][4]) || (phase_count[5] ^ phase[14][5]) || (phase_count[6] ^ phase[14][6]) || phase[14][7];
	assign select[15] = (phase_count[0] ^ phase[15][0]) || (phase_count[1] ^ phase[15][1]) || (phase_count[2] ^ phase[15][2]) || (phase_count[3] ^ phase[15][3]) || (phase_count[4] ^ phase[15][4]) || (phase_count[5] ^ phase[15][5]) || (phase_count[6] ^ phase[15][6]) || phase[15][7];
	assign select[16] = (phase_count[0] ^ phase[16][0]) || (phase_count[1] ^ phase[16][1]) || (phase_count[2] ^ phase[16][2]) || (phase_count[3] ^ phase[16][3]) || (phase_count[4] ^ phase[16][4]) || (phase_count[5] ^ phase[16][5]) || (phase_count[6] ^ phase[16][6]) || phase[16][7];
	assign select[17] = (phase_count[0] ^ phase[17][0]) || (phase_count[1] ^ phase[17][1]) || (phase_count[2] ^ phase[17][2]) || (phase_count[3] ^ phase[17][3]) || (phase_count[4] ^ phase[17][4]) || (phase_count[5] ^ phase[17][5]) || (phase_count[6] ^ phase[17][6]) || phase[17][7];
	assign select[18] = (phase_count[0] ^ phase[18][0]) || (phase_count[1] ^ phase[18][1]) || (phase_count[2] ^ phase[18][2]) || (phase_count[3] ^ phase[18][3]) || (phase_count[4] ^ phase[18][4]) || (phase_count[5] ^ phase[18][5]) || (phase_count[6] ^ phase[18][6]) || phase[18][7];
	assign select[19] = (phase_count[0] ^ phase[19][0]) || (phase_count[1] ^ phase[19][1]) || (phase_count[2] ^ phase[19][2]) || (phase_count[3] ^ phase[19][3]) || (phase_count[4] ^ phase[19][4]) || (phase_count[5] ^ phase[19][5]) || (phase_count[6] ^ phase[19][6]) || phase[19][7];
	assign select[20] = (phase_count[0] ^ phase[20][0]) || (phase_count[1] ^ phase[20][1]) || (phase_count[2] ^ phase[20][2]) || (phase_count[3] ^ phase[20][3]) || (phase_count[4] ^ phase[20][4]) || (phase_count[5] ^ phase[20][5]) || (phase_count[6] ^ phase[20][6]) || phase[20][7];
	assign select[21] = (phase_count[0] ^ phase[21][0]) || (phase_count[1] ^ phase[21][1]) || (phase_count[2] ^ phase[21][2]) || (phase_count[3] ^ phase[21][3]) || (phase_count[4] ^ phase[21][4]) || (phase_count[5] ^ phase[21][5]) || (phase_count[6] ^ phase[21][6]) || phase[21][7];
	assign select[22] = (phase_count[0] ^ phase[22][0]) || (phase_count[1] ^ phase[22][1]) || (phase_count[2] ^ phase[22][2]) || (phase_count[3] ^ phase[22][3]) || (phase_count[4] ^ phase[22][4]) || (phase_count[5] ^ phase[22][5]) || (phase_count[6] ^ phase[22][6]) || phase[22][7];
	assign select[23] = (phase_count[0] ^ phase[23][0]) || (phase_count[1] ^ phase[23][1]) || (phase_count[2] ^ phase[23][2]) || (phase_count[3] ^ phase[23][3]) || (phase_count[4] ^ phase[23][4]) || (phase_count[5] ^ phase[23][5]) || (phase_count[6] ^ phase[23][6]) || phase[23][7];
	assign select[24] = (phase_count[0] ^ phase[24][0]) || (phase_count[1] ^ phase[24][1]) || (phase_count[2] ^ phase[24][2]) || (phase_count[3] ^ phase[24][3]) || (phase_count[4] ^ phase[24][4]) || (phase_count[5] ^ phase[24][5]) || (phase_count[6] ^ phase[24][6]) || phase[24][7];
	assign select[25] = (phase_count[0] ^ phase[25][0]) || (phase_count[1] ^ phase[25][1]) || (phase_count[2] ^ phase[25][2]) || (phase_count[3] ^ phase[25][3]) || (phase_count[4] ^ phase[25][4]) || (phase_count[5] ^ phase[25][5]) || (phase_count[6] ^ phase[25][6]) || phase[25][7];
	assign select[26] = (phase_count[0] ^ phase[26][0]) || (phase_count[1] ^ phase[26][1]) || (phase_count[2] ^ phase[26][2]) || (phase_count[3] ^ phase[26][3]) || (phase_count[4] ^ phase[26][4]) || (phase_count[5] ^ phase[26][5]) || (phase_count[6] ^ phase[26][6]) || phase[26][7];
	assign select[27] = (phase_count[0] ^ phase[27][0]) || (phase_count[1] ^ phase[27][1]) || (phase_count[2] ^ phase[27][2]) || (phase_count[3] ^ phase[27][3]) || (phase_count[4] ^ phase[27][4]) || (phase_count[5] ^ phase[27][5]) || (phase_count[6] ^ phase[27][6]) || phase[27][7];
	assign select[28] = (phase_count[0] ^ phase[28][0]) || (phase_count[1] ^ phase[28][1]) || (phase_count[2] ^ phase[28][2]) || (phase_count[3] ^ phase[28][3]) || (phase_count[4] ^ phase[28][4]) || (phase_count[5] ^ phase[28][5]) || (phase_count[6] ^ phase[28][6]) || phase[28][7];
	assign select[29] = (phase_count[0] ^ phase[29][0]) || (phase_count[1] ^ phase[29][1]) || (phase_count[2] ^ phase[29][2]) || (phase_count[3] ^ phase[29][3]) || (phase_count[4] ^ phase[29][4]) || (phase_count[5] ^ phase[29][5]) || (phase_count[6] ^ phase[29][6]) || phase[29][7];
	assign select[30] = (phase_count[0] ^ phase[30][0]) || (phase_count[1] ^ phase[30][1]) || (phase_count[2] ^ phase[30][2]) || (phase_count[3] ^ phase[30][3]) || (phase_count[4] ^ phase[30][4]) || (phase_count[5] ^ phase[30][5]) || (phase_count[6] ^ phase[30][6]) || phase[30][7];
	assign select[31] = (phase_count[0] ^ phase[31][0]) || (phase_count[1] ^ phase[31][1]) || (phase_count[2] ^ phase[31][2]) || (phase_count[3] ^ phase[31][3]) || (phase_count[4] ^ phase[31][4]) || (phase_count[5] ^ phase[31][5]) || (phase_count[6] ^ phase[31][6]) || phase[31][7];
	assign select[32] = (phase_count[0] ^ phase[32][0]) || (phase_count[1] ^ phase[32][1]) || (phase_count[2] ^ phase[32][2]) || (phase_count[3] ^ phase[32][3]) || (phase_count[4] ^ phase[32][4]) || (phase_count[5] ^ phase[32][5]) || (phase_count[6] ^ phase[32][6]) || phase[32][7];
	assign select[33] = (phase_count[0] ^ phase[33][0]) || (phase_count[1] ^ phase[33][1]) || (phase_count[2] ^ phase[33][2]) || (phase_count[3] ^ phase[33][3]) || (phase_count[4] ^ phase[33][4]) || (phase_count[5] ^ phase[33][5]) || (phase_count[6] ^ phase[33][6]) || phase[33][7];
	assign select[34] = (phase_count[0] ^ phase[34][0]) || (phase_count[1] ^ phase[34][1]) || (phase_count[2] ^ phase[34][2]) || (phase_count[3] ^ phase[34][3]) || (phase_count[4] ^ phase[34][4]) || (phase_count[5] ^ phase[34][5]) || (phase_count[6] ^ phase[34][6]) || phase[34][7];
	assign select[35] = (phase_count[0] ^ phase[35][0]) || (phase_count[1] ^ phase[35][1]) || (phase_count[2] ^ phase[35][2]) || (phase_count[3] ^ phase[35][3]) || (phase_count[4] ^ phase[35][4]) || (phase_count[5] ^ phase[35][5]) || (phase_count[6] ^ phase[35][6]) || phase[35][7];
	assign select[36] = (phase_count[0] ^ phase[36][0]) || (phase_count[1] ^ phase[36][1]) || (phase_count[2] ^ phase[36][2]) || (phase_count[3] ^ phase[36][3]) || (phase_count[4] ^ phase[36][4]) || (phase_count[5] ^ phase[36][5]) || (phase_count[6] ^ phase[36][6]) || phase[36][7];
	assign select[37] = (phase_count[0] ^ phase[37][0]) || (phase_count[1] ^ phase[37][1]) || (phase_count[2] ^ phase[37][2]) || (phase_count[3] ^ phase[37][3]) || (phase_count[4] ^ phase[37][4]) || (phase_count[5] ^ phase[37][5]) || (phase_count[6] ^ phase[37][6]) || phase[37][7];
	assign select[38] = (phase_count[0] ^ phase[38][0]) || (phase_count[1] ^ phase[38][1]) || (phase_count[2] ^ phase[38][2]) || (phase_count[3] ^ phase[38][3]) || (phase_count[4] ^ phase[38][4]) || (phase_count[5] ^ phase[38][5]) || (phase_count[6] ^ phase[38][6]) || phase[38][7];
	assign select[39] = (phase_count[0] ^ phase[39][0]) || (phase_count[1] ^ phase[39][1]) || (phase_count[2] ^ phase[39][2]) || (phase_count[3] ^ phase[39][3]) || (phase_count[4] ^ phase[39][4]) || (phase_count[5] ^ phase[39][5]) || (phase_count[6] ^ phase[39][6]) || phase[39][7];
	assign select[40] = (phase_count[0] ^ phase[40][0]) || (phase_count[1] ^ phase[40][1]) || (phase_count[2] ^ phase[40][2]) || (phase_count[3] ^ phase[40][3]) || (phase_count[4] ^ phase[40][4]) || (phase_count[5] ^ phase[40][5]) || (phase_count[6] ^ phase[40][6]) || phase[40][7];
	assign select[41] = (phase_count[0] ^ phase[41][0]) || (phase_count[1] ^ phase[41][1]) || (phase_count[2] ^ phase[41][2]) || (phase_count[3] ^ phase[41][3]) || (phase_count[4] ^ phase[41][4]) || (phase_count[5] ^ phase[41][5]) || (phase_count[6] ^ phase[41][6]) || phase[41][7];
	assign select[42] = (phase_count[0] ^ phase[42][0]) || (phase_count[1] ^ phase[42][1]) || (phase_count[2] ^ phase[42][2]) || (phase_count[3] ^ phase[42][3]) || (phase_count[4] ^ phase[42][4]) || (phase_count[5] ^ phase[42][5]) || (phase_count[6] ^ phase[42][6]) || phase[42][7];
	assign select[43] = (phase_count[0] ^ phase[43][0]) || (phase_count[1] ^ phase[43][1]) || (phase_count[2] ^ phase[43][2]) || (phase_count[3] ^ phase[43][3]) || (phase_count[4] ^ phase[43][4]) || (phase_count[5] ^ phase[43][5]) || (phase_count[6] ^ phase[43][6]) || phase[43][7];
	assign select[44] = (phase_count[0] ^ phase[44][0]) || (phase_count[1] ^ phase[44][1]) || (phase_count[2] ^ phase[44][2]) || (phase_count[3] ^ phase[44][3]) || (phase_count[4] ^ phase[44][4]) || (phase_count[5] ^ phase[44][5]) || (phase_count[6] ^ phase[44][6]) || phase[44][7];
	assign select[45] = (phase_count[0] ^ phase[45][0]) || (phase_count[1] ^ phase[45][1]) || (phase_count[2] ^ phase[45][2]) || (phase_count[3] ^ phase[45][3]) || (phase_count[4] ^ phase[45][4]) || (phase_count[5] ^ phase[45][5]) || (phase_count[6] ^ phase[45][6]) || phase[45][7];
	assign select[46] = (phase_count[0] ^ phase[46][0]) || (phase_count[1] ^ phase[46][1]) || (phase_count[2] ^ phase[46][2]) || (phase_count[3] ^ phase[46][3]) || (phase_count[4] ^ phase[46][4]) || (phase_count[5] ^ phase[46][5]) || (phase_count[6] ^ phase[46][6]) || phase[46][7];
	assign select[47] = (phase_count[0] ^ phase[47][0]) || (phase_count[1] ^ phase[47][1]) || (phase_count[2] ^ phase[47][2]) || (phase_count[3] ^ phase[47][3]) || (phase_count[4] ^ phase[47][4]) || (phase_count[5] ^ phase[47][5]) || (phase_count[6] ^ phase[47][6]) || phase[47][7];
	assign select[48] = (phase_count[0] ^ phase[48][0]) || (phase_count[1] ^ phase[48][1]) || (phase_count[2] ^ phase[48][2]) || (phase_count[3] ^ phase[48][3]) || (phase_count[4] ^ phase[48][4]) || (phase_count[5] ^ phase[48][5]) || (phase_count[6] ^ phase[48][6]) || phase[48][7];
	assign select[49] = (phase_count[0] ^ phase[49][0]) || (phase_count[1] ^ phase[49][1]) || (phase_count[2] ^ phase[49][2]) || (phase_count[3] ^ phase[49][3]) || (phase_count[4] ^ phase[49][4]) || (phase_count[5] ^ phase[49][5]) || (phase_count[6] ^ phase[49][6]) || phase[49][7];
	assign select[50] = (phase_count[0] ^ phase[50][0]) || (phase_count[1] ^ phase[50][1]) || (phase_count[2] ^ phase[50][2]) || (phase_count[3] ^ phase[50][3]) || (phase_count[4] ^ phase[50][4]) || (phase_count[5] ^ phase[50][5]) || (phase_count[6] ^ phase[50][6]) || phase[50][7];
	assign select[51] = (phase_count[0] ^ phase[51][0]) || (phase_count[1] ^ phase[51][1]) || (phase_count[2] ^ phase[51][2]) || (phase_count[3] ^ phase[51][3]) || (phase_count[4] ^ phase[51][4]) || (phase_count[5] ^ phase[51][5]) || (phase_count[6] ^ phase[51][6]) || phase[51][7];
	assign select[52] = (phase_count[0] ^ phase[52][0]) || (phase_count[1] ^ phase[52][1]) || (phase_count[2] ^ phase[52][2]) || (phase_count[3] ^ phase[52][3]) || (phase_count[4] ^ phase[52][4]) || (phase_count[5] ^ phase[52][5]) || (phase_count[6] ^ phase[52][6]) || phase[52][7];
	assign select[53] = (phase_count[0] ^ phase[53][0]) || (phase_count[1] ^ phase[53][1]) || (phase_count[2] ^ phase[53][2]) || (phase_count[3] ^ phase[53][3]) || (phase_count[4] ^ phase[53][4]) || (phase_count[5] ^ phase[53][5]) || (phase_count[6] ^ phase[53][6]) || phase[53][7];
	assign select[54] = (phase_count[0] ^ phase[54][0]) || (phase_count[1] ^ phase[54][1]) || (phase_count[2] ^ phase[54][2]) || (phase_count[3] ^ phase[54][3]) || (phase_count[4] ^ phase[54][4]) || (phase_count[5] ^ phase[54][5]) || (phase_count[6] ^ phase[54][6]) || phase[54][7];
	assign select[55] = (phase_count[0] ^ phase[55][0]) || (phase_count[1] ^ phase[55][1]) || (phase_count[2] ^ phase[55][2]) || (phase_count[3] ^ phase[55][3]) || (phase_count[4] ^ phase[55][4]) || (phase_count[5] ^ phase[55][5]) || (phase_count[6] ^ phase[55][6]) || phase[55][7];
	assign select[56] = (phase_count[0] ^ phase[56][0]) || (phase_count[1] ^ phase[56][1]) || (phase_count[2] ^ phase[56][2]) || (phase_count[3] ^ phase[56][3]) || (phase_count[4] ^ phase[56][4]) || (phase_count[5] ^ phase[56][5]) || (phase_count[6] ^ phase[56][6]) || phase[56][7];
	assign select[57] = (phase_count[0] ^ phase[57][0]) || (phase_count[1] ^ phase[57][1]) || (phase_count[2] ^ phase[57][2]) || (phase_count[3] ^ phase[57][3]) || (phase_count[4] ^ phase[57][4]) || (phase_count[5] ^ phase[57][5]) || (phase_count[6] ^ phase[57][6]) || phase[57][7];
	assign select[58] = (phase_count[0] ^ phase[58][0]) || (phase_count[1] ^ phase[58][1]) || (phase_count[2] ^ phase[58][2]) || (phase_count[3] ^ phase[58][3]) || (phase_count[4] ^ phase[58][4]) || (phase_count[5] ^ phase[58][5]) || (phase_count[6] ^ phase[58][6]) || phase[58][7];
	assign select[59] = (phase_count[0] ^ phase[59][0]) || (phase_count[1] ^ phase[59][1]) || (phase_count[2] ^ phase[59][2]) || (phase_count[3] ^ phase[59][3]) || (phase_count[4] ^ phase[59][4]) || (phase_count[5] ^ phase[59][5]) || (phase_count[6] ^ phase[59][6]) || phase[59][7];
	assign select[60] = (phase_count[0] ^ phase[60][0]) || (phase_count[1] ^ phase[60][1]) || (phase_count[2] ^ phase[60][2]) || (phase_count[3] ^ phase[60][3]) || (phase_count[4] ^ phase[60][4]) || (phase_count[5] ^ phase[60][5]) || (phase_count[6] ^ phase[60][6]) || phase[60][7];
	assign select[61] = (phase_count[0] ^ phase[61][0]) || (phase_count[1] ^ phase[61][1]) || (phase_count[2] ^ phase[61][2]) || (phase_count[3] ^ phase[61][3]) || (phase_count[4] ^ phase[61][4]) || (phase_count[5] ^ phase[61][5]) || (phase_count[6] ^ phase[61][6]) || phase[61][7];
	assign select[62] = (phase_count[0] ^ phase[62][0]) || (phase_count[1] ^ phase[62][1]) || (phase_count[2] ^ phase[62][2]) || (phase_count[3] ^ phase[62][3]) || (phase_count[4] ^ phase[62][4]) || (phase_count[5] ^ phase[62][5]) || (phase_count[6] ^ phase[62][6]) || phase[62][7];
	assign select[63] = (phase_count[0] ^ phase[63][0]) || (phase_count[1] ^ phase[63][1]) || (phase_count[2] ^ phase[63][2]) || (phase_count[3] ^ phase[63][3]) || (phase_count[4] ^ phase[63][4]) || (phase_count[5] ^ phase[63][5]) || (phase_count[6] ^ phase[63][6]) || phase[63][7];
	assign select[64] = (phase_count[0] ^ phase[64][0]) || (phase_count[1] ^ phase[64][1]) || (phase_count[2] ^ phase[64][2]) || (phase_count[3] ^ phase[64][3]) || (phase_count[4] ^ phase[64][4]) || (phase_count[5] ^ phase[64][5]) || (phase_count[6] ^ phase[64][6]) || phase[64][7];
	assign select[65] = (phase_count[0] ^ phase[65][0]) || (phase_count[1] ^ phase[65][1]) || (phase_count[2] ^ phase[65][2]) || (phase_count[3] ^ phase[65][3]) || (phase_count[4] ^ phase[65][4]) || (phase_count[5] ^ phase[65][5]) || (phase_count[6] ^ phase[65][6]) || phase[65][7];
	assign select[66] = (phase_count[0] ^ phase[66][0]) || (phase_count[1] ^ phase[66][1]) || (phase_count[2] ^ phase[66][2]) || (phase_count[3] ^ phase[66][3]) || (phase_count[4] ^ phase[66][4]) || (phase_count[5] ^ phase[66][5]) || (phase_count[6] ^ phase[66][6]) || phase[66][7];
	assign select[67] = (phase_count[0] ^ phase[67][0]) || (phase_count[1] ^ phase[67][1]) || (phase_count[2] ^ phase[67][2]) || (phase_count[3] ^ phase[67][3]) || (phase_count[4] ^ phase[67][4]) || (phase_count[5] ^ phase[67][5]) || (phase_count[6] ^ phase[67][6]) || phase[67][7];
	assign select[68] = (phase_count[0] ^ phase[68][0]) || (phase_count[1] ^ phase[68][1]) || (phase_count[2] ^ phase[68][2]) || (phase_count[3] ^ phase[68][3]) || (phase_count[4] ^ phase[68][4]) || (phase_count[5] ^ phase[68][5]) || (phase_count[6] ^ phase[68][6]) || phase[68][7];
	assign select[69] = (phase_count[0] ^ phase[69][0]) || (phase_count[1] ^ phase[69][1]) || (phase_count[2] ^ phase[69][2]) || (phase_count[3] ^ phase[69][3]) || (phase_count[4] ^ phase[69][4]) || (phase_count[5] ^ phase[69][5]) || (phase_count[6] ^ phase[69][6]) || phase[69][7];
	assign select[70] = (phase_count[0] ^ phase[70][0]) || (phase_count[1] ^ phase[70][1]) || (phase_count[2] ^ phase[70][2]) || (phase_count[3] ^ phase[70][3]) || (phase_count[4] ^ phase[70][4]) || (phase_count[5] ^ phase[70][5]) || (phase_count[6] ^ phase[70][6]) || phase[70][7];
	assign select[71] = (phase_count[0] ^ phase[71][0]) || (phase_count[1] ^ phase[71][1]) || (phase_count[2] ^ phase[71][2]) || (phase_count[3] ^ phase[71][3]) || (phase_count[4] ^ phase[71][4]) || (phase_count[5] ^ phase[71][5]) || (phase_count[6] ^ phase[71][6]) || phase[71][7];
	assign select[72] = (phase_count[0] ^ phase[72][0]) || (phase_count[1] ^ phase[72][1]) || (phase_count[2] ^ phase[72][2]) || (phase_count[3] ^ phase[72][3]) || (phase_count[4] ^ phase[72][4]) || (phase_count[5] ^ phase[72][5]) || (phase_count[6] ^ phase[72][6]) || phase[72][7];
	assign select[73] = (phase_count[0] ^ phase[73][0]) || (phase_count[1] ^ phase[73][1]) || (phase_count[2] ^ phase[73][2]) || (phase_count[3] ^ phase[73][3]) || (phase_count[4] ^ phase[73][4]) || (phase_count[5] ^ phase[73][5]) || (phase_count[6] ^ phase[73][6]) || phase[73][7];
	assign select[74] = (phase_count[0] ^ phase[74][0]) || (phase_count[1] ^ phase[74][1]) || (phase_count[2] ^ phase[74][2]) || (phase_count[3] ^ phase[74][3]) || (phase_count[4] ^ phase[74][4]) || (phase_count[5] ^ phase[74][5]) || (phase_count[6] ^ phase[74][6]) || phase[74][7];
	assign select[75] = (phase_count[0] ^ phase[75][0]) || (phase_count[1] ^ phase[75][1]) || (phase_count[2] ^ phase[75][2]) || (phase_count[3] ^ phase[75][3]) || (phase_count[4] ^ phase[75][4]) || (phase_count[5] ^ phase[75][5]) || (phase_count[6] ^ phase[75][6]) || phase[75][7];
	assign select[76] = (phase_count[0] ^ phase[76][0]) || (phase_count[1] ^ phase[76][1]) || (phase_count[2] ^ phase[76][2]) || (phase_count[3] ^ phase[76][3]) || (phase_count[4] ^ phase[76][4]) || (phase_count[5] ^ phase[76][5]) || (phase_count[6] ^ phase[76][6]) || phase[76][7];
	assign select[77] = (phase_count[0] ^ phase[77][0]) || (phase_count[1] ^ phase[77][1]) || (phase_count[2] ^ phase[77][2]) || (phase_count[3] ^ phase[77][3]) || (phase_count[4] ^ phase[77][4]) || (phase_count[5] ^ phase[77][5]) || (phase_count[6] ^ phase[77][6]) || phase[77][7];
	assign select[78] = (phase_count[0] ^ phase[78][0]) || (phase_count[1] ^ phase[78][1]) || (phase_count[2] ^ phase[78][2]) || (phase_count[3] ^ phase[78][3]) || (phase_count[4] ^ phase[78][4]) || (phase_count[5] ^ phase[78][5]) || (phase_count[6] ^ phase[78][6]) || phase[78][7];
	assign select[79] = (phase_count[0] ^ phase[79][0]) || (phase_count[1] ^ phase[79][1]) || (phase_count[2] ^ phase[79][2]) || (phase_count[3] ^ phase[79][3]) || (phase_count[4] ^ phase[79][4]) || (phase_count[5] ^ phase[79][5]) || (phase_count[6] ^ phase[79][6]) || phase[79][7];
	assign select[80] = (phase_count[0] ^ phase[80][0]) || (phase_count[1] ^ phase[80][1]) || (phase_count[2] ^ phase[80][2]) || (phase_count[3] ^ phase[80][3]) || (phase_count[4] ^ phase[80][4]) || (phase_count[5] ^ phase[80][5]) || (phase_count[6] ^ phase[80][6]) || phase[80][7];
	assign select[81] = (phase_count[0] ^ phase[81][0]) || (phase_count[1] ^ phase[81][1]) || (phase_count[2] ^ phase[81][2]) || (phase_count[3] ^ phase[81][3]) || (phase_count[4] ^ phase[81][4]) || (phase_count[5] ^ phase[81][5]) || (phase_count[6] ^ phase[81][6]) || phase[81][7];
	assign select[82] = (phase_count[0] ^ phase[82][0]) || (phase_count[1] ^ phase[82][1]) || (phase_count[2] ^ phase[82][2]) || (phase_count[3] ^ phase[82][3]) || (phase_count[4] ^ phase[82][4]) || (phase_count[5] ^ phase[82][5]) || (phase_count[6] ^ phase[82][6]) || phase[82][7];
	assign select[83] = (phase_count[0] ^ phase[83][0]) || (phase_count[1] ^ phase[83][1]) || (phase_count[2] ^ phase[83][2]) || (phase_count[3] ^ phase[83][3]) || (phase_count[4] ^ phase[83][4]) || (phase_count[5] ^ phase[83][5]) || (phase_count[6] ^ phase[83][6]) || phase[83][7];
	assign select[84] = (phase_count[0] ^ phase[84][0]) || (phase_count[1] ^ phase[84][1]) || (phase_count[2] ^ phase[84][2]) || (phase_count[3] ^ phase[84][3]) || (phase_count[4] ^ phase[84][4]) || (phase_count[5] ^ phase[84][5]) || (phase_count[6] ^ phase[84][6]) || phase[84][7];
	assign select[85] = (phase_count[0] ^ phase[85][0]) || (phase_count[1] ^ phase[85][1]) || (phase_count[2] ^ phase[85][2]) || (phase_count[3] ^ phase[85][3]) || (phase_count[4] ^ phase[85][4]) || (phase_count[5] ^ phase[85][5]) || (phase_count[6] ^ phase[85][6]) || phase[85][7];
	assign select[86] = (phase_count[0] ^ phase[86][0]) || (phase_count[1] ^ phase[86][1]) || (phase_count[2] ^ phase[86][2]) || (phase_count[3] ^ phase[86][3]) || (phase_count[4] ^ phase[86][4]) || (phase_count[5] ^ phase[86][5]) || (phase_count[6] ^ phase[86][6]) || phase[86][7];
	assign select[87] = (phase_count[0] ^ phase[87][0]) || (phase_count[1] ^ phase[87][1]) || (phase_count[2] ^ phase[87][2]) || (phase_count[3] ^ phase[87][3]) || (phase_count[4] ^ phase[87][4]) || (phase_count[5] ^ phase[87][5]) || (phase_count[6] ^ phase[87][6]) || phase[87][7];
	assign select[88] = (phase_count[0] ^ phase[88][0]) || (phase_count[1] ^ phase[88][1]) || (phase_count[2] ^ phase[88][2]) || (phase_count[3] ^ phase[88][3]) || (phase_count[4] ^ phase[88][4]) || (phase_count[5] ^ phase[88][5]) || (phase_count[6] ^ phase[88][6]) || phase[88][7];
	assign select[89] = (phase_count[0] ^ phase[89][0]) || (phase_count[1] ^ phase[89][1]) || (phase_count[2] ^ phase[89][2]) || (phase_count[3] ^ phase[89][3]) || (phase_count[4] ^ phase[89][4]) || (phase_count[5] ^ phase[89][5]) || (phase_count[6] ^ phase[89][6]) || phase[89][7];
	assign select[90] = (phase_count[0] ^ phase[90][0]) || (phase_count[1] ^ phase[90][1]) || (phase_count[2] ^ phase[90][2]) || (phase_count[3] ^ phase[90][3]) || (phase_count[4] ^ phase[90][4]) || (phase_count[5] ^ phase[90][5]) || (phase_count[6] ^ phase[90][6]) || phase[90][7];
	assign select[91] = (phase_count[0] ^ phase[91][0]) || (phase_count[1] ^ phase[91][1]) || (phase_count[2] ^ phase[91][2]) || (phase_count[3] ^ phase[91][3]) || (phase_count[4] ^ phase[91][4]) || (phase_count[5] ^ phase[91][5]) || (phase_count[6] ^ phase[91][6]) || phase[91][7];
	assign select[92] = (phase_count[0] ^ phase[92][0]) || (phase_count[1] ^ phase[92][1]) || (phase_count[2] ^ phase[92][2]) || (phase_count[3] ^ phase[92][3]) || (phase_count[4] ^ phase[92][4]) || (phase_count[5] ^ phase[92][5]) || (phase_count[6] ^ phase[92][6]) || phase[92][7];
	assign select[93] = (phase_count[0] ^ phase[93][0]) || (phase_count[1] ^ phase[93][1]) || (phase_count[2] ^ phase[93][2]) || (phase_count[3] ^ phase[93][3]) || (phase_count[4] ^ phase[93][4]) || (phase_count[5] ^ phase[93][5]) || (phase_count[6] ^ phase[93][6]) || phase[93][7];
	assign select[94] = (phase_count[0] ^ phase[94][0]) || (phase_count[1] ^ phase[94][1]) || (phase_count[2] ^ phase[94][2]) || (phase_count[3] ^ phase[94][3]) || (phase_count[4] ^ phase[94][4]) || (phase_count[5] ^ phase[94][5]) || (phase_count[6] ^ phase[94][6]) || phase[94][7];
	assign select[95] = (phase_count[0] ^ phase[95][0]) || (phase_count[1] ^ phase[95][1]) || (phase_count[2] ^ phase[95][2]) || (phase_count[3] ^ phase[95][3]) || (phase_count[4] ^ phase[95][4]) || (phase_count[5] ^ phase[95][5]) || (phase_count[6] ^ phase[95][6]) || phase[95][7];
	assign select[96] = (phase_count[0] ^ phase[96][0]) || (phase_count[1] ^ phase[96][1]) || (phase_count[2] ^ phase[96][2]) || (phase_count[3] ^ phase[96][3]) || (phase_count[4] ^ phase[96][4]) || (phase_count[5] ^ phase[96][5]) || (phase_count[6] ^ phase[96][6]) || phase[96][7];
	assign select[97] = (phase_count[0] ^ phase[97][0]) || (phase_count[1] ^ phase[97][1]) || (phase_count[2] ^ phase[97][2]) || (phase_count[3] ^ phase[97][3]) || (phase_count[4] ^ phase[97][4]) || (phase_count[5] ^ phase[97][5]) || (phase_count[6] ^ phase[97][6]) || phase[97][7];
	assign select[98] = (phase_count[0] ^ phase[98][0]) || (phase_count[1] ^ phase[98][1]) || (phase_count[2] ^ phase[98][2]) || (phase_count[3] ^ phase[98][3]) || (phase_count[4] ^ phase[98][4]) || (phase_count[5] ^ phase[98][5]) || (phase_count[6] ^ phase[98][6]) || phase[98][7];
	assign select[99] = (phase_count[0] ^ phase[99][0]) || (phase_count[1] ^ phase[99][1]) || (phase_count[2] ^ phase[99][2]) || (phase_count[3] ^ phase[99][3]) || (phase_count[4] ^ phase[99][4]) || (phase_count[5] ^ phase[99][5]) || (phase_count[6] ^ phase[99][6]) || phase[99][7];
	assign select[100] = (phase_count[0] ^ phase[100][0]) || (phase_count[1] ^ phase[100][1]) || (phase_count[2] ^ phase[100][2]) || (phase_count[3] ^ phase[100][3]) || (phase_count[4] ^ phase[100][4]) || (phase_count[5] ^ phase[100][5]) || (phase_count[6] ^ phase[100][6]) || phase[100][7];
	assign select[101] = (phase_count[0] ^ phase[101][0]) || (phase_count[1] ^ phase[101][1]) || (phase_count[2] ^ phase[101][2]) || (phase_count[3] ^ phase[101][3]) || (phase_count[4] ^ phase[101][4]) || (phase_count[5] ^ phase[101][5]) || (phase_count[6] ^ phase[101][6]) || phase[101][7];
	assign select[102] = (phase_count[0] ^ phase[102][0]) || (phase_count[1] ^ phase[102][1]) || (phase_count[2] ^ phase[102][2]) || (phase_count[3] ^ phase[102][3]) || (phase_count[4] ^ phase[102][4]) || (phase_count[5] ^ phase[102][5]) || (phase_count[6] ^ phase[102][6]) || phase[102][7];
	assign select[103] = (phase_count[0] ^ phase[103][0]) || (phase_count[1] ^ phase[103][1]) || (phase_count[2] ^ phase[103][2]) || (phase_count[3] ^ phase[103][3]) || (phase_count[4] ^ phase[103][4]) || (phase_count[5] ^ phase[103][5]) || (phase_count[6] ^ phase[103][6]) || phase[103][7];
	assign select[104] = (phase_count[0] ^ phase[104][0]) || (phase_count[1] ^ phase[104][1]) || (phase_count[2] ^ phase[104][2]) || (phase_count[3] ^ phase[104][3]) || (phase_count[4] ^ phase[104][4]) || (phase_count[5] ^ phase[104][5]) || (phase_count[6] ^ phase[104][6]) || phase[104][7];
	assign select[105] = (phase_count[0] ^ phase[105][0]) || (phase_count[1] ^ phase[105][1]) || (phase_count[2] ^ phase[105][2]) || (phase_count[3] ^ phase[105][3]) || (phase_count[4] ^ phase[105][4]) || (phase_count[5] ^ phase[105][5]) || (phase_count[6] ^ phase[105][6]) || phase[105][7];
	assign select[106] = (phase_count[0] ^ phase[106][0]) || (phase_count[1] ^ phase[106][1]) || (phase_count[2] ^ phase[106][2]) || (phase_count[3] ^ phase[106][3]) || (phase_count[4] ^ phase[106][4]) || (phase_count[5] ^ phase[106][5]) || (phase_count[6] ^ phase[106][6]) || phase[106][7];
	assign select[107] = (phase_count[0] ^ phase[107][0]) || (phase_count[1] ^ phase[107][1]) || (phase_count[2] ^ phase[107][2]) || (phase_count[3] ^ phase[107][3]) || (phase_count[4] ^ phase[107][4]) || (phase_count[5] ^ phase[107][5]) || (phase_count[6] ^ phase[107][6]) || phase[107][7];
	assign select[108] = (phase_count[0] ^ phase[108][0]) || (phase_count[1] ^ phase[108][1]) || (phase_count[2] ^ phase[108][2]) || (phase_count[3] ^ phase[108][3]) || (phase_count[4] ^ phase[108][4]) || (phase_count[5] ^ phase[108][5]) || (phase_count[6] ^ phase[108][6]) || phase[108][7];
	assign select[109] = (phase_count[0] ^ phase[109][0]) || (phase_count[1] ^ phase[109][1]) || (phase_count[2] ^ phase[109][2]) || (phase_count[3] ^ phase[109][3]) || (phase_count[4] ^ phase[109][4]) || (phase_count[5] ^ phase[109][5]) || (phase_count[6] ^ phase[109][6]) || phase[109][7];
	assign select[110] = (phase_count[0] ^ phase[110][0]) || (phase_count[1] ^ phase[110][1]) || (phase_count[2] ^ phase[110][2]) || (phase_count[3] ^ phase[110][3]) || (phase_count[4] ^ phase[110][4]) || (phase_count[5] ^ phase[110][5]) || (phase_count[6] ^ phase[110][6]) || phase[110][7];
	assign select[111] = (phase_count[0] ^ phase[111][0]) || (phase_count[1] ^ phase[111][1]) || (phase_count[2] ^ phase[111][2]) || (phase_count[3] ^ phase[111][3]) || (phase_count[4] ^ phase[111][4]) || (phase_count[5] ^ phase[111][5]) || (phase_count[6] ^ phase[111][6]) || phase[111][7];
	assign select[112] = (phase_count[0] ^ phase[112][0]) || (phase_count[1] ^ phase[112][1]) || (phase_count[2] ^ phase[112][2]) || (phase_count[3] ^ phase[112][3]) || (phase_count[4] ^ phase[112][4]) || (phase_count[5] ^ phase[112][5]) || (phase_count[6] ^ phase[112][6]) || phase[112][7];
	assign select[113] = (phase_count[0] ^ phase[113][0]) || (phase_count[1] ^ phase[113][1]) || (phase_count[2] ^ phase[113][2]) || (phase_count[3] ^ phase[113][3]) || (phase_count[4] ^ phase[113][4]) || (phase_count[5] ^ phase[113][5]) || (phase_count[6] ^ phase[113][6]) || phase[113][7];
	assign select[114] = (phase_count[0] ^ phase[114][0]) || (phase_count[1] ^ phase[114][1]) || (phase_count[2] ^ phase[114][2]) || (phase_count[3] ^ phase[114][3]) || (phase_count[4] ^ phase[114][4]) || (phase_count[5] ^ phase[114][5]) || (phase_count[6] ^ phase[114][6]) || phase[114][7];
	assign select[115] = (phase_count[0] ^ phase[115][0]) || (phase_count[1] ^ phase[115][1]) || (phase_count[2] ^ phase[115][2]) || (phase_count[3] ^ phase[115][3]) || (phase_count[4] ^ phase[115][4]) || (phase_count[5] ^ phase[115][5]) || (phase_count[6] ^ phase[115][6]) || phase[115][7];
	assign select[116] = (phase_count[0] ^ phase[116][0]) || (phase_count[1] ^ phase[116][1]) || (phase_count[2] ^ phase[116][2]) || (phase_count[3] ^ phase[116][3]) || (phase_count[4] ^ phase[116][4]) || (phase_count[5] ^ phase[116][5]) || (phase_count[6] ^ phase[116][6]) || phase[116][7];
	assign select[117] = (phase_count[0] ^ phase[117][0]) || (phase_count[1] ^ phase[117][1]) || (phase_count[2] ^ phase[117][2]) || (phase_count[3] ^ phase[117][3]) || (phase_count[4] ^ phase[117][4]) || (phase_count[5] ^ phase[117][5]) || (phase_count[6] ^ phase[117][6]) || phase[117][7];
	assign select[118] = (phase_count[0] ^ phase[118][0]) || (phase_count[1] ^ phase[118][1]) || (phase_count[2] ^ phase[118][2]) || (phase_count[3] ^ phase[118][3]) || (phase_count[4] ^ phase[118][4]) || (phase_count[5] ^ phase[118][5]) || (phase_count[6] ^ phase[118][6]) || phase[118][7];
	assign select[119] = (phase_count[0] ^ phase[119][0]) || (phase_count[1] ^ phase[119][1]) || (phase_count[2] ^ phase[119][2]) || (phase_count[3] ^ phase[119][3]) || (phase_count[4] ^ phase[119][4]) || (phase_count[5] ^ phase[119][5]) || (phase_count[6] ^ phase[119][6]) || phase[119][7];
	assign select[120] = (phase_count[0] ^ phase[120][0]) || (phase_count[1] ^ phase[120][1]) || (phase_count[2] ^ phase[120][2]) || (phase_count[3] ^ phase[120][3]) || (phase_count[4] ^ phase[120][4]) || (phase_count[5] ^ phase[120][5]) || (phase_count[6] ^ phase[120][6]) || phase[120][7];
	assign select[121] = (phase_count[0] ^ phase[121][0]) || (phase_count[1] ^ phase[121][1]) || (phase_count[2] ^ phase[121][2]) || (phase_count[3] ^ phase[121][3]) || (phase_count[4] ^ phase[121][4]) || (phase_count[5] ^ phase[121][5]) || (phase_count[6] ^ phase[121][6]) || phase[121][7];
	assign select[122] = (phase_count[0] ^ phase[122][0]) || (phase_count[1] ^ phase[122][1]) || (phase_count[2] ^ phase[122][2]) || (phase_count[3] ^ phase[122][3]) || (phase_count[4] ^ phase[122][4]) || (phase_count[5] ^ phase[122][5]) || (phase_count[6] ^ phase[122][6]) || phase[122][7];
	assign select[123] = (phase_count[0] ^ phase[123][0]) || (phase_count[1] ^ phase[123][1]) || (phase_count[2] ^ phase[123][2]) || (phase_count[3] ^ phase[123][3]) || (phase_count[4] ^ phase[123][4]) || (phase_count[5] ^ phase[123][5]) || (phase_count[6] ^ phase[123][6]) || phase[123][7];
	assign select[124] = (phase_count[0] ^ phase[124][0]) || (phase_count[1] ^ phase[124][1]) || (phase_count[2] ^ phase[124][2]) || (phase_count[3] ^ phase[124][3]) || (phase_count[4] ^ phase[124][4]) || (phase_count[5] ^ phase[124][5]) || (phase_count[6] ^ phase[124][6]) || phase[124][7];
	assign select[125] = (phase_count[0] ^ phase[125][0]) || (phase_count[1] ^ phase[125][1]) || (phase_count[2] ^ phase[125][2]) || (phase_count[3] ^ phase[125][3]) || (phase_count[4] ^ phase[125][4]) || (phase_count[5] ^ phase[125][5]) || (phase_count[6] ^ phase[125][6]) || phase[125][7];
	assign select[126] = (phase_count[0] ^ phase[126][0]) || (phase_count[1] ^ phase[126][1]) || (phase_count[2] ^ phase[126][2]) || (phase_count[3] ^ phase[126][3]) || (phase_count[4] ^ phase[126][4]) || (phase_count[5] ^ phase[126][5]) || (phase_count[6] ^ phase[126][6]) || phase[126][7];
	assign select[127] = (phase_count[0] ^ phase[127][0]) || (phase_count[1] ^ phase[127][1]) || (phase_count[2] ^ phase[127][2]) || (phase_count[3] ^ phase[127][3]) || (phase_count[4] ^ phase[127][4]) || (phase_count[5] ^ phase[127][5]) || (phase_count[6] ^ phase[127][6]) || phase[127][7];
	assign select[128] = (phase_count[0] ^ phase[128][0]) || (phase_count[1] ^ phase[128][1]) || (phase_count[2] ^ phase[128][2]) || (phase_count[3] ^ phase[128][3]) || (phase_count[4] ^ phase[128][4]) || (phase_count[5] ^ phase[128][5]) || (phase_count[6] ^ phase[128][6]) || phase[128][7];
	assign select[129] = (phase_count[0] ^ phase[129][0]) || (phase_count[1] ^ phase[129][1]) || (phase_count[2] ^ phase[129][2]) || (phase_count[3] ^ phase[129][3]) || (phase_count[4] ^ phase[129][4]) || (phase_count[5] ^ phase[129][5]) || (phase_count[6] ^ phase[129][6]) || phase[129][7];
	assign select[130] = (phase_count[0] ^ phase[130][0]) || (phase_count[1] ^ phase[130][1]) || (phase_count[2] ^ phase[130][2]) || (phase_count[3] ^ phase[130][3]) || (phase_count[4] ^ phase[130][4]) || (phase_count[5] ^ phase[130][5]) || (phase_count[6] ^ phase[130][6]) || phase[130][7];
	assign select[131] = (phase_count[0] ^ phase[131][0]) || (phase_count[1] ^ phase[131][1]) || (phase_count[2] ^ phase[131][2]) || (phase_count[3] ^ phase[131][3]) || (phase_count[4] ^ phase[131][4]) || (phase_count[5] ^ phase[131][5]) || (phase_count[6] ^ phase[131][6]) || phase[131][7];
	assign select[132] = (phase_count[0] ^ phase[132][0]) || (phase_count[1] ^ phase[132][1]) || (phase_count[2] ^ phase[132][2]) || (phase_count[3] ^ phase[132][3]) || (phase_count[4] ^ phase[132][4]) || (phase_count[5] ^ phase[132][5]) || (phase_count[6] ^ phase[132][6]) || phase[132][7];
	assign select[133] = (phase_count[0] ^ phase[133][0]) || (phase_count[1] ^ phase[133][1]) || (phase_count[2] ^ phase[133][2]) || (phase_count[3] ^ phase[133][3]) || (phase_count[4] ^ phase[133][4]) || (phase_count[5] ^ phase[133][5]) || (phase_count[6] ^ phase[133][6]) || phase[133][7];
	assign select[134] = (phase_count[0] ^ phase[134][0]) || (phase_count[1] ^ phase[134][1]) || (phase_count[2] ^ phase[134][2]) || (phase_count[3] ^ phase[134][3]) || (phase_count[4] ^ phase[134][4]) || (phase_count[5] ^ phase[134][5]) || (phase_count[6] ^ phase[134][6]) || phase[134][7];
	assign select[135] = (phase_count[0] ^ phase[135][0]) || (phase_count[1] ^ phase[135][1]) || (phase_count[2] ^ phase[135][2]) || (phase_count[3] ^ phase[135][3]) || (phase_count[4] ^ phase[135][4]) || (phase_count[5] ^ phase[135][5]) || (phase_count[6] ^ phase[135][6]) || phase[135][7];
	assign select[136] = (phase_count[0] ^ phase[136][0]) || (phase_count[1] ^ phase[136][1]) || (phase_count[2] ^ phase[136][2]) || (phase_count[3] ^ phase[136][3]) || (phase_count[4] ^ phase[136][4]) || (phase_count[5] ^ phase[136][5]) || (phase_count[6] ^ phase[136][6]) || phase[136][7];
	assign select[137] = (phase_count[0] ^ phase[137][0]) || (phase_count[1] ^ phase[137][1]) || (phase_count[2] ^ phase[137][2]) || (phase_count[3] ^ phase[137][3]) || (phase_count[4] ^ phase[137][4]) || (phase_count[5] ^ phase[137][5]) || (phase_count[6] ^ phase[137][6]) || phase[137][7];
	assign select[138] = (phase_count[0] ^ phase[138][0]) || (phase_count[1] ^ phase[138][1]) || (phase_count[2] ^ phase[138][2]) || (phase_count[3] ^ phase[138][3]) || (phase_count[4] ^ phase[138][4]) || (phase_count[5] ^ phase[138][5]) || (phase_count[6] ^ phase[138][6]) || phase[138][7];
	assign select[139] = (phase_count[0] ^ phase[139][0]) || (phase_count[1] ^ phase[139][1]) || (phase_count[2] ^ phase[139][2]) || (phase_count[3] ^ phase[139][3]) || (phase_count[4] ^ phase[139][4]) || (phase_count[5] ^ phase[139][5]) || (phase_count[6] ^ phase[139][6]) || phase[139][7];
	assign select[140] = (phase_count[0] ^ phase[140][0]) || (phase_count[1] ^ phase[140][1]) || (phase_count[2] ^ phase[140][2]) || (phase_count[3] ^ phase[140][3]) || (phase_count[4] ^ phase[140][4]) || (phase_count[5] ^ phase[140][5]) || (phase_count[6] ^ phase[140][6]) || phase[140][7];
	assign select[141] = (phase_count[0] ^ phase[141][0]) || (phase_count[1] ^ phase[141][1]) || (phase_count[2] ^ phase[141][2]) || (phase_count[3] ^ phase[141][3]) || (phase_count[4] ^ phase[141][4]) || (phase_count[5] ^ phase[141][5]) || (phase_count[6] ^ phase[141][6]) || phase[141][7];
	assign select[142] = (phase_count[0] ^ phase[142][0]) || (phase_count[1] ^ phase[142][1]) || (phase_count[2] ^ phase[142][2]) || (phase_count[3] ^ phase[142][3]) || (phase_count[4] ^ phase[142][4]) || (phase_count[5] ^ phase[142][5]) || (phase_count[6] ^ phase[142][6]) || phase[142][7];
	assign select[143] = (phase_count[0] ^ phase[143][0]) || (phase_count[1] ^ phase[143][1]) || (phase_count[2] ^ phase[143][2]) || (phase_count[3] ^ phase[143][3]) || (phase_count[4] ^ phase[143][4]) || (phase_count[5] ^ phase[143][5]) || (phase_count[6] ^ phase[143][6]) || phase[143][7];
	assign select[144] = (phase_count[0] ^ phase[144][0]) || (phase_count[1] ^ phase[144][1]) || (phase_count[2] ^ phase[144][2]) || (phase_count[3] ^ phase[144][3]) || (phase_count[4] ^ phase[144][4]) || (phase_count[5] ^ phase[144][5]) || (phase_count[6] ^ phase[144][6]) || phase[144][7];
	assign select[145] = (phase_count[0] ^ phase[145][0]) || (phase_count[1] ^ phase[145][1]) || (phase_count[2] ^ phase[145][2]) || (phase_count[3] ^ phase[145][3]) || (phase_count[4] ^ phase[145][4]) || (phase_count[5] ^ phase[145][5]) || (phase_count[6] ^ phase[145][6]) || phase[145][7];
	assign select[146] = (phase_count[0] ^ phase[146][0]) || (phase_count[1] ^ phase[146][1]) || (phase_count[2] ^ phase[146][2]) || (phase_count[3] ^ phase[146][3]) || (phase_count[4] ^ phase[146][4]) || (phase_count[5] ^ phase[146][5]) || (phase_count[6] ^ phase[146][6]) || phase[146][7];
	assign select[147] = (phase_count[0] ^ phase[147][0]) || (phase_count[1] ^ phase[147][1]) || (phase_count[2] ^ phase[147][2]) || (phase_count[3] ^ phase[147][3]) || (phase_count[4] ^ phase[147][4]) || (phase_count[5] ^ phase[147][5]) || (phase_count[6] ^ phase[147][6]) || phase[147][7];
	assign select[148] = (phase_count[0] ^ phase[148][0]) || (phase_count[1] ^ phase[148][1]) || (phase_count[2] ^ phase[148][2]) || (phase_count[3] ^ phase[148][3]) || (phase_count[4] ^ phase[148][4]) || (phase_count[5] ^ phase[148][5]) || (phase_count[6] ^ phase[148][6]) || phase[148][7];
	assign select[149] = (phase_count[0] ^ phase[149][0]) || (phase_count[1] ^ phase[149][1]) || (phase_count[2] ^ phase[149][2]) || (phase_count[3] ^ phase[149][3]) || (phase_count[4] ^ phase[149][4]) || (phase_count[5] ^ phase[149][5]) || (phase_count[6] ^ phase[149][6]) || phase[149][7];
	assign select[150] = (phase_count[0] ^ phase[150][0]) || (phase_count[1] ^ phase[150][1]) || (phase_count[2] ^ phase[150][2]) || (phase_count[3] ^ phase[150][3]) || (phase_count[4] ^ phase[150][4]) || (phase_count[5] ^ phase[150][5]) || (phase_count[6] ^ phase[150][6]) || phase[150][7];
	assign select[151] = (phase_count[0] ^ phase[151][0]) || (phase_count[1] ^ phase[151][1]) || (phase_count[2] ^ phase[151][2]) || (phase_count[3] ^ phase[151][3]) || (phase_count[4] ^ phase[151][4]) || (phase_count[5] ^ phase[151][5]) || (phase_count[6] ^ phase[151][6]) || phase[151][7];
	assign select[152] = (phase_count[0] ^ phase[152][0]) || (phase_count[1] ^ phase[152][1]) || (phase_count[2] ^ phase[152][2]) || (phase_count[3] ^ phase[152][3]) || (phase_count[4] ^ phase[152][4]) || (phase_count[5] ^ phase[152][5]) || (phase_count[6] ^ phase[152][6]) || phase[152][7];
	assign select[153] = (phase_count[0] ^ phase[153][0]) || (phase_count[1] ^ phase[153][1]) || (phase_count[2] ^ phase[153][2]) || (phase_count[3] ^ phase[153][3]) || (phase_count[4] ^ phase[153][4]) || (phase_count[5] ^ phase[153][5]) || (phase_count[6] ^ phase[153][6]) || phase[153][7];
	assign select[154] = (phase_count[0] ^ phase[154][0]) || (phase_count[1] ^ phase[154][1]) || (phase_count[2] ^ phase[154][2]) || (phase_count[3] ^ phase[154][3]) || (phase_count[4] ^ phase[154][4]) || (phase_count[5] ^ phase[154][5]) || (phase_count[6] ^ phase[154][6]) || phase[154][7];
	assign select[155] = (phase_count[0] ^ phase[155][0]) || (phase_count[1] ^ phase[155][1]) || (phase_count[2] ^ phase[155][2]) || (phase_count[3] ^ phase[155][3]) || (phase_count[4] ^ phase[155][4]) || (phase_count[5] ^ phase[155][5]) || (phase_count[6] ^ phase[155][6]) || phase[155][7];
	assign select[156] = (phase_count[0] ^ phase[156][0]) || (phase_count[1] ^ phase[156][1]) || (phase_count[2] ^ phase[156][2]) || (phase_count[3] ^ phase[156][3]) || (phase_count[4] ^ phase[156][4]) || (phase_count[5] ^ phase[156][5]) || (phase_count[6] ^ phase[156][6]) || phase[156][7];
	assign select[157] = (phase_count[0] ^ phase[157][0]) || (phase_count[1] ^ phase[157][1]) || (phase_count[2] ^ phase[157][2]) || (phase_count[3] ^ phase[157][3]) || (phase_count[4] ^ phase[157][4]) || (phase_count[5] ^ phase[157][5]) || (phase_count[6] ^ phase[157][6]) || phase[157][7];
	assign select[158] = (phase_count[0] ^ phase[158][0]) || (phase_count[1] ^ phase[158][1]) || (phase_count[2] ^ phase[158][2]) || (phase_count[3] ^ phase[158][3]) || (phase_count[4] ^ phase[158][4]) || (phase_count[5] ^ phase[158][5]) || (phase_count[6] ^ phase[158][6]) || phase[158][7];
	assign select[159] = (phase_count[0] ^ phase[159][0]) || (phase_count[1] ^ phase[159][1]) || (phase_count[2] ^ phase[159][2]) || (phase_count[3] ^ phase[159][3]) || (phase_count[4] ^ phase[159][4]) || (phase_count[5] ^ phase[159][5]) || (phase_count[6] ^ phase[159][6]) || phase[159][7];
	assign select[160] = (phase_count[0] ^ phase[160][0]) || (phase_count[1] ^ phase[160][1]) || (phase_count[2] ^ phase[160][2]) || (phase_count[3] ^ phase[160][3]) || (phase_count[4] ^ phase[160][4]) || (phase_count[5] ^ phase[160][5]) || (phase_count[6] ^ phase[160][6]) || phase[160][7];
	assign select[161] = (phase_count[0] ^ phase[161][0]) || (phase_count[1] ^ phase[161][1]) || (phase_count[2] ^ phase[161][2]) || (phase_count[3] ^ phase[161][3]) || (phase_count[4] ^ phase[161][4]) || (phase_count[5] ^ phase[161][5]) || (phase_count[6] ^ phase[161][6]) || phase[161][7];
	assign select[162] = (phase_count[0] ^ phase[162][0]) || (phase_count[1] ^ phase[162][1]) || (phase_count[2] ^ phase[162][2]) || (phase_count[3] ^ phase[162][3]) || (phase_count[4] ^ phase[162][4]) || (phase_count[5] ^ phase[162][5]) || (phase_count[6] ^ phase[162][6]) || phase[162][7];
	assign select[163] = (phase_count[0] ^ phase[163][0]) || (phase_count[1] ^ phase[163][1]) || (phase_count[2] ^ phase[163][2]) || (phase_count[3] ^ phase[163][3]) || (phase_count[4] ^ phase[163][4]) || (phase_count[5] ^ phase[163][5]) || (phase_count[6] ^ phase[163][6]) || phase[163][7];
	assign select[164] = (phase_count[0] ^ phase[164][0]) || (phase_count[1] ^ phase[164][1]) || (phase_count[2] ^ phase[164][2]) || (phase_count[3] ^ phase[164][3]) || (phase_count[4] ^ phase[164][4]) || (phase_count[5] ^ phase[164][5]) || (phase_count[6] ^ phase[164][6]) || phase[164][7];
	assign select[165] = (phase_count[0] ^ phase[165][0]) || (phase_count[1] ^ phase[165][1]) || (phase_count[2] ^ phase[165][2]) || (phase_count[3] ^ phase[165][3]) || (phase_count[4] ^ phase[165][4]) || (phase_count[5] ^ phase[165][5]) || (phase_count[6] ^ phase[165][6]) || phase[165][7];
	assign select[166] = (phase_count[0] ^ phase[166][0]) || (phase_count[1] ^ phase[166][1]) || (phase_count[2] ^ phase[166][2]) || (phase_count[3] ^ phase[166][3]) || (phase_count[4] ^ phase[166][4]) || (phase_count[5] ^ phase[166][5]) || (phase_count[6] ^ phase[166][6]) || phase[166][7];
	assign select[167] = (phase_count[0] ^ phase[167][0]) || (phase_count[1] ^ phase[167][1]) || (phase_count[2] ^ phase[167][2]) || (phase_count[3] ^ phase[167][3]) || (phase_count[4] ^ phase[167][4]) || (phase_count[5] ^ phase[167][5]) || (phase_count[6] ^ phase[167][6]) || phase[167][7];
	assign select[168] = (phase_count[0] ^ phase[168][0]) || (phase_count[1] ^ phase[168][1]) || (phase_count[2] ^ phase[168][2]) || (phase_count[3] ^ phase[168][3]) || (phase_count[4] ^ phase[168][4]) || (phase_count[5] ^ phase[168][5]) || (phase_count[6] ^ phase[168][6]) || phase[168][7];
	assign select[169] = (phase_count[0] ^ phase[169][0]) || (phase_count[1] ^ phase[169][1]) || (phase_count[2] ^ phase[169][2]) || (phase_count[3] ^ phase[169][3]) || (phase_count[4] ^ phase[169][4]) || (phase_count[5] ^ phase[169][5]) || (phase_count[6] ^ phase[169][6]) || phase[169][7];
	assign select[170] = (phase_count[0] ^ phase[170][0]) || (phase_count[1] ^ phase[170][1]) || (phase_count[2] ^ phase[170][2]) || (phase_count[3] ^ phase[170][3]) || (phase_count[4] ^ phase[170][4]) || (phase_count[5] ^ phase[170][5]) || (phase_count[6] ^ phase[170][6]) || phase[170][7];
	assign select[171] = (phase_count[0] ^ phase[171][0]) || (phase_count[1] ^ phase[171][1]) || (phase_count[2] ^ phase[171][2]) || (phase_count[3] ^ phase[171][3]) || (phase_count[4] ^ phase[171][4]) || (phase_count[5] ^ phase[171][5]) || (phase_count[6] ^ phase[171][6]) || phase[171][7];
	assign select[172] = (phase_count[0] ^ phase[172][0]) || (phase_count[1] ^ phase[172][1]) || (phase_count[2] ^ phase[172][2]) || (phase_count[3] ^ phase[172][3]) || (phase_count[4] ^ phase[172][4]) || (phase_count[5] ^ phase[172][5]) || (phase_count[6] ^ phase[172][6]) || phase[172][7];
	assign select[173] = (phase_count[0] ^ phase[173][0]) || (phase_count[1] ^ phase[173][1]) || (phase_count[2] ^ phase[173][2]) || (phase_count[3] ^ phase[173][3]) || (phase_count[4] ^ phase[173][4]) || (phase_count[5] ^ phase[173][5]) || (phase_count[6] ^ phase[173][6]) || phase[173][7];
	assign select[174] = (phase_count[0] ^ phase[174][0]) || (phase_count[1] ^ phase[174][1]) || (phase_count[2] ^ phase[174][2]) || (phase_count[3] ^ phase[174][3]) || (phase_count[4] ^ phase[174][4]) || (phase_count[5] ^ phase[174][5]) || (phase_count[6] ^ phase[174][6]) || phase[174][7];
	assign select[175] = (phase_count[0] ^ phase[175][0]) || (phase_count[1] ^ phase[175][1]) || (phase_count[2] ^ phase[175][2]) || (phase_count[3] ^ phase[175][3]) || (phase_count[4] ^ phase[175][4]) || (phase_count[5] ^ phase[175][5]) || (phase_count[6] ^ phase[175][6]) || phase[175][7];
	assign select[176] = (phase_count[0] ^ phase[176][0]) || (phase_count[1] ^ phase[176][1]) || (phase_count[2] ^ phase[176][2]) || (phase_count[3] ^ phase[176][3]) || (phase_count[4] ^ phase[176][4]) || (phase_count[5] ^ phase[176][5]) || (phase_count[6] ^ phase[176][6]) || phase[176][7];
	assign select[177] = (phase_count[0] ^ phase[177][0]) || (phase_count[1] ^ phase[177][1]) || (phase_count[2] ^ phase[177][2]) || (phase_count[3] ^ phase[177][3]) || (phase_count[4] ^ phase[177][4]) || (phase_count[5] ^ phase[177][5]) || (phase_count[6] ^ phase[177][6]) || phase[177][7];
	assign select[178] = (phase_count[0] ^ phase[178][0]) || (phase_count[1] ^ phase[178][1]) || (phase_count[2] ^ phase[178][2]) || (phase_count[3] ^ phase[178][3]) || (phase_count[4] ^ phase[178][4]) || (phase_count[5] ^ phase[178][5]) || (phase_count[6] ^ phase[178][6]) || phase[178][7];
	assign select[179] = (phase_count[0] ^ phase[179][0]) || (phase_count[1] ^ phase[179][1]) || (phase_count[2] ^ phase[179][2]) || (phase_count[3] ^ phase[179][3]) || (phase_count[4] ^ phase[179][4]) || (phase_count[5] ^ phase[179][5]) || (phase_count[6] ^ phase[179][6]) || phase[179][7];
	assign select[180] = (phase_count[0] ^ phase[180][0]) || (phase_count[1] ^ phase[180][1]) || (phase_count[2] ^ phase[180][2]) || (phase_count[3] ^ phase[180][3]) || (phase_count[4] ^ phase[180][4]) || (phase_count[5] ^ phase[180][5]) || (phase_count[6] ^ phase[180][6]) || phase[180][7];
	assign select[181] = (phase_count[0] ^ phase[181][0]) || (phase_count[1] ^ phase[181][1]) || (phase_count[2] ^ phase[181][2]) || (phase_count[3] ^ phase[181][3]) || (phase_count[4] ^ phase[181][4]) || (phase_count[5] ^ phase[181][5]) || (phase_count[6] ^ phase[181][6]) || phase[181][7];
	assign select[182] = (phase_count[0] ^ phase[182][0]) || (phase_count[1] ^ phase[182][1]) || (phase_count[2] ^ phase[182][2]) || (phase_count[3] ^ phase[182][3]) || (phase_count[4] ^ phase[182][4]) || (phase_count[5] ^ phase[182][5]) || (phase_count[6] ^ phase[182][6]) || phase[182][7];
	assign select[183] = (phase_count[0] ^ phase[183][0]) || (phase_count[1] ^ phase[183][1]) || (phase_count[2] ^ phase[183][2]) || (phase_count[3] ^ phase[183][3]) || (phase_count[4] ^ phase[183][4]) || (phase_count[5] ^ phase[183][5]) || (phase_count[6] ^ phase[183][6]) || phase[183][7];
	assign select[184] = (phase_count[0] ^ phase[184][0]) || (phase_count[1] ^ phase[184][1]) || (phase_count[2] ^ phase[184][2]) || (phase_count[3] ^ phase[184][3]) || (phase_count[4] ^ phase[184][4]) || (phase_count[5] ^ phase[184][5]) || (phase_count[6] ^ phase[184][6]) || phase[184][7];
	assign select[185] = (phase_count[0] ^ phase[185][0]) || (phase_count[1] ^ phase[185][1]) || (phase_count[2] ^ phase[185][2]) || (phase_count[3] ^ phase[185][3]) || (phase_count[4] ^ phase[185][4]) || (phase_count[5] ^ phase[185][5]) || (phase_count[6] ^ phase[185][6]) || phase[185][7];
	assign select[186] = (phase_count[0] ^ phase[186][0]) || (phase_count[1] ^ phase[186][1]) || (phase_count[2] ^ phase[186][2]) || (phase_count[3] ^ phase[186][3]) || (phase_count[4] ^ phase[186][4]) || (phase_count[5] ^ phase[186][5]) || (phase_count[6] ^ phase[186][6]) || phase[186][7];
	assign select[187] = (phase_count[0] ^ phase[187][0]) || (phase_count[1] ^ phase[187][1]) || (phase_count[2] ^ phase[187][2]) || (phase_count[3] ^ phase[187][3]) || (phase_count[4] ^ phase[187][4]) || (phase_count[5] ^ phase[187][5]) || (phase_count[6] ^ phase[187][6]) || phase[187][7];
	assign select[188] = (phase_count[0] ^ phase[188][0]) || (phase_count[1] ^ phase[188][1]) || (phase_count[2] ^ phase[188][2]) || (phase_count[3] ^ phase[188][3]) || (phase_count[4] ^ phase[188][4]) || (phase_count[5] ^ phase[188][5]) || (phase_count[6] ^ phase[188][6]) || phase[188][7];
	assign select[189] = (phase_count[0] ^ phase[189][0]) || (phase_count[1] ^ phase[189][1]) || (phase_count[2] ^ phase[189][2]) || (phase_count[3] ^ phase[189][3]) || (phase_count[4] ^ phase[189][4]) || (phase_count[5] ^ phase[189][5]) || (phase_count[6] ^ phase[189][6]) || phase[189][7];
	assign select[190] = (phase_count[0] ^ phase[190][0]) || (phase_count[1] ^ phase[190][1]) || (phase_count[2] ^ phase[190][2]) || (phase_count[3] ^ phase[190][3]) || (phase_count[4] ^ phase[190][4]) || (phase_count[5] ^ phase[190][5]) || (phase_count[6] ^ phase[190][6]) || phase[190][7];
	assign select[191] = (phase_count[0] ^ phase[191][0]) || (phase_count[1] ^ phase[191][1]) || (phase_count[2] ^ phase[191][2]) || (phase_count[3] ^ phase[191][3]) || (phase_count[4] ^ phase[191][4]) || (phase_count[5] ^ phase[191][5]) || (phase_count[6] ^ phase[191][6]) || phase[191][7];
	assign select[192] = (phase_count[0] ^ phase[192][0]) || (phase_count[1] ^ phase[192][1]) || (phase_count[2] ^ phase[192][2]) || (phase_count[3] ^ phase[192][3]) || (phase_count[4] ^ phase[192][4]) || (phase_count[5] ^ phase[192][5]) || (phase_count[6] ^ phase[192][6]) || phase[192][7];
	assign select[193] = (phase_count[0] ^ phase[193][0]) || (phase_count[1] ^ phase[193][1]) || (phase_count[2] ^ phase[193][2]) || (phase_count[3] ^ phase[193][3]) || (phase_count[4] ^ phase[193][4]) || (phase_count[5] ^ phase[193][5]) || (phase_count[6] ^ phase[193][6]) || phase[193][7];
	assign select[194] = (phase_count[0] ^ phase[194][0]) || (phase_count[1] ^ phase[194][1]) || (phase_count[2] ^ phase[194][2]) || (phase_count[3] ^ phase[194][3]) || (phase_count[4] ^ phase[194][4]) || (phase_count[5] ^ phase[194][5]) || (phase_count[6] ^ phase[194][6]) || phase[194][7];
	assign select[195] = (phase_count[0] ^ phase[195][0]) || (phase_count[1] ^ phase[195][1]) || (phase_count[2] ^ phase[195][2]) || (phase_count[3] ^ phase[195][3]) || (phase_count[4] ^ phase[195][4]) || (phase_count[5] ^ phase[195][5]) || (phase_count[6] ^ phase[195][6]) || phase[195][7];
	assign select[196] = (phase_count[0] ^ phase[196][0]) || (phase_count[1] ^ phase[196][1]) || (phase_count[2] ^ phase[196][2]) || (phase_count[3] ^ phase[196][3]) || (phase_count[4] ^ phase[196][4]) || (phase_count[5] ^ phase[196][5]) || (phase_count[6] ^ phase[196][6]) || phase[196][7];
	assign select[197] = (phase_count[0] ^ phase[197][0]) || (phase_count[1] ^ phase[197][1]) || (phase_count[2] ^ phase[197][2]) || (phase_count[3] ^ phase[197][3]) || (phase_count[4] ^ phase[197][4]) || (phase_count[5] ^ phase[197][5]) || (phase_count[6] ^ phase[197][6]) || phase[197][7];
	assign select[198] = (phase_count[0] ^ phase[198][0]) || (phase_count[1] ^ phase[198][1]) || (phase_count[2] ^ phase[198][2]) || (phase_count[3] ^ phase[198][3]) || (phase_count[4] ^ phase[198][4]) || (phase_count[5] ^ phase[198][5]) || (phase_count[6] ^ phase[198][6]) || phase[198][7];
	assign select[199] = (phase_count[0] ^ phase[199][0]) || (phase_count[1] ^ phase[199][1]) || (phase_count[2] ^ phase[199][2]) || (phase_count[3] ^ phase[199][3]) || (phase_count[4] ^ phase[199][4]) || (phase_count[5] ^ phase[199][5]) || (phase_count[6] ^ phase[199][6]) || phase[199][7];
	assign select[200] = (phase_count[0] ^ phase[200][0]) || (phase_count[1] ^ phase[200][1]) || (phase_count[2] ^ phase[200][2]) || (phase_count[3] ^ phase[200][3]) || (phase_count[4] ^ phase[200][4]) || (phase_count[5] ^ phase[200][5]) || (phase_count[6] ^ phase[200][6]) || phase[200][7];
	assign select[201] = (phase_count[0] ^ phase[201][0]) || (phase_count[1] ^ phase[201][1]) || (phase_count[2] ^ phase[201][2]) || (phase_count[3] ^ phase[201][3]) || (phase_count[4] ^ phase[201][4]) || (phase_count[5] ^ phase[201][5]) || (phase_count[6] ^ phase[201][6]) || phase[201][7];
	assign select[202] = (phase_count[0] ^ phase[202][0]) || (phase_count[1] ^ phase[202][1]) || (phase_count[2] ^ phase[202][2]) || (phase_count[3] ^ phase[202][3]) || (phase_count[4] ^ phase[202][4]) || (phase_count[5] ^ phase[202][5]) || (phase_count[6] ^ phase[202][6]) || phase[202][7];
	assign select[203] = (phase_count[0] ^ phase[203][0]) || (phase_count[1] ^ phase[203][1]) || (phase_count[2] ^ phase[203][2]) || (phase_count[3] ^ phase[203][3]) || (phase_count[4] ^ phase[203][4]) || (phase_count[5] ^ phase[203][5]) || (phase_count[6] ^ phase[203][6]) || phase[203][7];
	assign select[204] = (phase_count[0] ^ phase[204][0]) || (phase_count[1] ^ phase[204][1]) || (phase_count[2] ^ phase[204][2]) || (phase_count[3] ^ phase[204][3]) || (phase_count[4] ^ phase[204][4]) || (phase_count[5] ^ phase[204][5]) || (phase_count[6] ^ phase[204][6]) || phase[204][7];
	assign select[205] = (phase_count[0] ^ phase[205][0]) || (phase_count[1] ^ phase[205][1]) || (phase_count[2] ^ phase[205][2]) || (phase_count[3] ^ phase[205][3]) || (phase_count[4] ^ phase[205][4]) || (phase_count[5] ^ phase[205][5]) || (phase_count[6] ^ phase[205][6]) || phase[205][7];
	assign select[206] = (phase_count[0] ^ phase[206][0]) || (phase_count[1] ^ phase[206][1]) || (phase_count[2] ^ phase[206][2]) || (phase_count[3] ^ phase[206][3]) || (phase_count[4] ^ phase[206][4]) || (phase_count[5] ^ phase[206][5]) || (phase_count[6] ^ phase[206][6]) || phase[206][7];
	assign select[207] = (phase_count[0] ^ phase[207][0]) || (phase_count[1] ^ phase[207][1]) || (phase_count[2] ^ phase[207][2]) || (phase_count[3] ^ phase[207][3]) || (phase_count[4] ^ phase[207][4]) || (phase_count[5] ^ phase[207][5]) || (phase_count[6] ^ phase[207][6]) || phase[207][7];
	assign select[208] = (phase_count[0] ^ phase[208][0]) || (phase_count[1] ^ phase[208][1]) || (phase_count[2] ^ phase[208][2]) || (phase_count[3] ^ phase[208][3]) || (phase_count[4] ^ phase[208][4]) || (phase_count[5] ^ phase[208][5]) || (phase_count[6] ^ phase[208][6]) || phase[208][7];
	assign select[209] = (phase_count[0] ^ phase[209][0]) || (phase_count[1] ^ phase[209][1]) || (phase_count[2] ^ phase[209][2]) || (phase_count[3] ^ phase[209][3]) || (phase_count[4] ^ phase[209][4]) || (phase_count[5] ^ phase[209][5]) || (phase_count[6] ^ phase[209][6]) || phase[209][7];
	assign select[210] = (phase_count[0] ^ phase[210][0]) || (phase_count[1] ^ phase[210][1]) || (phase_count[2] ^ phase[210][2]) || (phase_count[3] ^ phase[210][3]) || (phase_count[4] ^ phase[210][4]) || (phase_count[5] ^ phase[210][5]) || (phase_count[6] ^ phase[210][6]) || phase[210][7];
	assign select[211] = (phase_count[0] ^ phase[211][0]) || (phase_count[1] ^ phase[211][1]) || (phase_count[2] ^ phase[211][2]) || (phase_count[3] ^ phase[211][3]) || (phase_count[4] ^ phase[211][4]) || (phase_count[5] ^ phase[211][5]) || (phase_count[6] ^ phase[211][6]) || phase[211][7];
	assign select[212] = (phase_count[0] ^ phase[212][0]) || (phase_count[1] ^ phase[212][1]) || (phase_count[2] ^ phase[212][2]) || (phase_count[3] ^ phase[212][3]) || (phase_count[4] ^ phase[212][4]) || (phase_count[5] ^ phase[212][5]) || (phase_count[6] ^ phase[212][6]) || phase[212][7];
	assign select[213] = (phase_count[0] ^ phase[213][0]) || (phase_count[1] ^ phase[213][1]) || (phase_count[2] ^ phase[213][2]) || (phase_count[3] ^ phase[213][3]) || (phase_count[4] ^ phase[213][4]) || (phase_count[5] ^ phase[213][5]) || (phase_count[6] ^ phase[213][6]) || phase[213][7];
	assign select[214] = (phase_count[0] ^ phase[214][0]) || (phase_count[1] ^ phase[214][1]) || (phase_count[2] ^ phase[214][2]) || (phase_count[3] ^ phase[214][3]) || (phase_count[4] ^ phase[214][4]) || (phase_count[5] ^ phase[214][5]) || (phase_count[6] ^ phase[214][6]) || phase[214][7];
	assign select[215] = (phase_count[0] ^ phase[215][0]) || (phase_count[1] ^ phase[215][1]) || (phase_count[2] ^ phase[215][2]) || (phase_count[3] ^ phase[215][3]) || (phase_count[4] ^ phase[215][4]) || (phase_count[5] ^ phase[215][5]) || (phase_count[6] ^ phase[215][6]) || phase[215][7];
	assign select[216] = (phase_count[0] ^ phase[216][0]) || (phase_count[1] ^ phase[216][1]) || (phase_count[2] ^ phase[216][2]) || (phase_count[3] ^ phase[216][3]) || (phase_count[4] ^ phase[216][4]) || (phase_count[5] ^ phase[216][5]) || (phase_count[6] ^ phase[216][6]) || phase[216][7];
	assign select[217] = (phase_count[0] ^ phase[217][0]) || (phase_count[1] ^ phase[217][1]) || (phase_count[2] ^ phase[217][2]) || (phase_count[3] ^ phase[217][3]) || (phase_count[4] ^ phase[217][4]) || (phase_count[5] ^ phase[217][5]) || (phase_count[6] ^ phase[217][6]) || phase[217][7];
	assign select[218] = (phase_count[0] ^ phase[218][0]) || (phase_count[1] ^ phase[218][1]) || (phase_count[2] ^ phase[218][2]) || (phase_count[3] ^ phase[218][3]) || (phase_count[4] ^ phase[218][4]) || (phase_count[5] ^ phase[218][5]) || (phase_count[6] ^ phase[218][6]) || phase[218][7];
	assign select[219] = (phase_count[0] ^ phase[219][0]) || (phase_count[1] ^ phase[219][1]) || (phase_count[2] ^ phase[219][2]) || (phase_count[3] ^ phase[219][3]) || (phase_count[4] ^ phase[219][4]) || (phase_count[5] ^ phase[219][5]) || (phase_count[6] ^ phase[219][6]) || phase[219][7];
	assign select[220] = (phase_count[0] ^ phase[220][0]) || (phase_count[1] ^ phase[220][1]) || (phase_count[2] ^ phase[220][2]) || (phase_count[3] ^ phase[220][3]) || (phase_count[4] ^ phase[220][4]) || (phase_count[5] ^ phase[220][5]) || (phase_count[6] ^ phase[220][6]) || phase[220][7];
	assign select[221] = (phase_count[0] ^ phase[221][0]) || (phase_count[1] ^ phase[221][1]) || (phase_count[2] ^ phase[221][2]) || (phase_count[3] ^ phase[221][3]) || (phase_count[4] ^ phase[221][4]) || (phase_count[5] ^ phase[221][5]) || (phase_count[6] ^ phase[221][6]) || phase[221][7];
	assign select[222] = (phase_count[0] ^ phase[222][0]) || (phase_count[1] ^ phase[222][1]) || (phase_count[2] ^ phase[222][2]) || (phase_count[3] ^ phase[222][3]) || (phase_count[4] ^ phase[222][4]) || (phase_count[5] ^ phase[222][5]) || (phase_count[6] ^ phase[222][6]) || phase[222][7];
	assign select[223] = (phase_count[0] ^ phase[223][0]) || (phase_count[1] ^ phase[223][1]) || (phase_count[2] ^ phase[223][2]) || (phase_count[3] ^ phase[223][3]) || (phase_count[4] ^ phase[223][4]) || (phase_count[5] ^ phase[223][5]) || (phase_count[6] ^ phase[223][6]) || phase[223][7];
	assign select[224] = (phase_count[0] ^ phase[224][0]) || (phase_count[1] ^ phase[224][1]) || (phase_count[2] ^ phase[224][2]) || (phase_count[3] ^ phase[224][3]) || (phase_count[4] ^ phase[224][4]) || (phase_count[5] ^ phase[224][5]) || (phase_count[6] ^ phase[224][6]) || phase[224][7];
	assign select[225] = (phase_count[0] ^ phase[225][0]) || (phase_count[1] ^ phase[225][1]) || (phase_count[2] ^ phase[225][2]) || (phase_count[3] ^ phase[225][3]) || (phase_count[4] ^ phase[225][4]) || (phase_count[5] ^ phase[225][5]) || (phase_count[6] ^ phase[225][6]) || phase[225][7];
	assign select[226] = (phase_count[0] ^ phase[226][0]) || (phase_count[1] ^ phase[226][1]) || (phase_count[2] ^ phase[226][2]) || (phase_count[3] ^ phase[226][3]) || (phase_count[4] ^ phase[226][4]) || (phase_count[5] ^ phase[226][5]) || (phase_count[6] ^ phase[226][6]) || phase[226][7];
	assign select[227] = (phase_count[0] ^ phase[227][0]) || (phase_count[1] ^ phase[227][1]) || (phase_count[2] ^ phase[227][2]) || (phase_count[3] ^ phase[227][3]) || (phase_count[4] ^ phase[227][4]) || (phase_count[5] ^ phase[227][5]) || (phase_count[6] ^ phase[227][6]) || phase[227][7];
	assign select[228] = (phase_count[0] ^ phase[228][0]) || (phase_count[1] ^ phase[228][1]) || (phase_count[2] ^ phase[228][2]) || (phase_count[3] ^ phase[228][3]) || (phase_count[4] ^ phase[228][4]) || (phase_count[5] ^ phase[228][5]) || (phase_count[6] ^ phase[228][6]) || phase[228][7];
	assign select[229] = (phase_count[0] ^ phase[229][0]) || (phase_count[1] ^ phase[229][1]) || (phase_count[2] ^ phase[229][2]) || (phase_count[3] ^ phase[229][3]) || (phase_count[4] ^ phase[229][4]) || (phase_count[5] ^ phase[229][5]) || (phase_count[6] ^ phase[229][6]) || phase[229][7];
	assign select[230] = (phase_count[0] ^ phase[230][0]) || (phase_count[1] ^ phase[230][1]) || (phase_count[2] ^ phase[230][2]) || (phase_count[3] ^ phase[230][3]) || (phase_count[4] ^ phase[230][4]) || (phase_count[5] ^ phase[230][5]) || (phase_count[6] ^ phase[230][6]) || phase[230][7];
	assign select[231] = (phase_count[0] ^ phase[231][0]) || (phase_count[1] ^ phase[231][1]) || (phase_count[2] ^ phase[231][2]) || (phase_count[3] ^ phase[231][3]) || (phase_count[4] ^ phase[231][4]) || (phase_count[5] ^ phase[231][5]) || (phase_count[6] ^ phase[231][6]) || phase[231][7];
	assign select[232] = (phase_count[0] ^ phase[232][0]) || (phase_count[1] ^ phase[232][1]) || (phase_count[2] ^ phase[232][2]) || (phase_count[3] ^ phase[232][3]) || (phase_count[4] ^ phase[232][4]) || (phase_count[5] ^ phase[232][5]) || (phase_count[6] ^ phase[232][6]) || phase[232][7];
	assign select[233] = (phase_count[0] ^ phase[233][0]) || (phase_count[1] ^ phase[233][1]) || (phase_count[2] ^ phase[233][2]) || (phase_count[3] ^ phase[233][3]) || (phase_count[4] ^ phase[233][4]) || (phase_count[5] ^ phase[233][5]) || (phase_count[6] ^ phase[233][6]) || phase[233][7];
	assign select[234] = (phase_count[0] ^ phase[234][0]) || (phase_count[1] ^ phase[234][1]) || (phase_count[2] ^ phase[234][2]) || (phase_count[3] ^ phase[234][3]) || (phase_count[4] ^ phase[234][4]) || (phase_count[5] ^ phase[234][5]) || (phase_count[6] ^ phase[234][6]) || phase[234][7];
	assign select[235] = (phase_count[0] ^ phase[235][0]) || (phase_count[1] ^ phase[235][1]) || (phase_count[2] ^ phase[235][2]) || (phase_count[3] ^ phase[235][3]) || (phase_count[4] ^ phase[235][4]) || (phase_count[5] ^ phase[235][5]) || (phase_count[6] ^ phase[235][6]) || phase[235][7];
	assign select[236] = (phase_count[0] ^ phase[236][0]) || (phase_count[1] ^ phase[236][1]) || (phase_count[2] ^ phase[236][2]) || (phase_count[3] ^ phase[236][3]) || (phase_count[4] ^ phase[236][4]) || (phase_count[5] ^ phase[236][5]) || (phase_count[6] ^ phase[236][6]) || phase[236][7];
	assign select[237] = (phase_count[0] ^ phase[237][0]) || (phase_count[1] ^ phase[237][1]) || (phase_count[2] ^ phase[237][2]) || (phase_count[3] ^ phase[237][3]) || (phase_count[4] ^ phase[237][4]) || (phase_count[5] ^ phase[237][5]) || (phase_count[6] ^ phase[237][6]) || phase[237][7];
	assign select[238] = (phase_count[0] ^ phase[238][0]) || (phase_count[1] ^ phase[238][1]) || (phase_count[2] ^ phase[238][2]) || (phase_count[3] ^ phase[238][3]) || (phase_count[4] ^ phase[238][4]) || (phase_count[5] ^ phase[238][5]) || (phase_count[6] ^ phase[238][6]) || phase[238][7];
	assign select[239] = (phase_count[0] ^ phase[239][0]) || (phase_count[1] ^ phase[239][1]) || (phase_count[2] ^ phase[239][2]) || (phase_count[3] ^ phase[239][3]) || (phase_count[4] ^ phase[239][4]) || (phase_count[5] ^ phase[239][5]) || (phase_count[6] ^ phase[239][6]) || phase[239][7];
	assign select[240] = (phase_count[0] ^ phase[240][0]) || (phase_count[1] ^ phase[240][1]) || (phase_count[2] ^ phase[240][2]) || (phase_count[3] ^ phase[240][3]) || (phase_count[4] ^ phase[240][4]) || (phase_count[5] ^ phase[240][5]) || (phase_count[6] ^ phase[240][6]) || phase[240][7];
	assign select[241] = (phase_count[0] ^ phase[241][0]) || (phase_count[1] ^ phase[241][1]) || (phase_count[2] ^ phase[241][2]) || (phase_count[3] ^ phase[241][3]) || (phase_count[4] ^ phase[241][4]) || (phase_count[5] ^ phase[241][5]) || (phase_count[6] ^ phase[241][6]) || phase[241][7];
	assign select[242] = (phase_count[0] ^ phase[242][0]) || (phase_count[1] ^ phase[242][1]) || (phase_count[2] ^ phase[242][2]) || (phase_count[3] ^ phase[242][3]) || (phase_count[4] ^ phase[242][4]) || (phase_count[5] ^ phase[242][5]) || (phase_count[6] ^ phase[242][6]) || phase[242][7];
	assign select[243] = (phase_count[0] ^ phase[243][0]) || (phase_count[1] ^ phase[243][1]) || (phase_count[2] ^ phase[243][2]) || (phase_count[3] ^ phase[243][3]) || (phase_count[4] ^ phase[243][4]) || (phase_count[5] ^ phase[243][5]) || (phase_count[6] ^ phase[243][6]) || phase[243][7];
	assign select[244] = (phase_count[0] ^ phase[244][0]) || (phase_count[1] ^ phase[244][1]) || (phase_count[2] ^ phase[244][2]) || (phase_count[3] ^ phase[244][3]) || (phase_count[4] ^ phase[244][4]) || (phase_count[5] ^ phase[244][5]) || (phase_count[6] ^ phase[244][6]) || phase[244][7];
	assign select[245] = (phase_count[0] ^ phase[245][0]) || (phase_count[1] ^ phase[245][1]) || (phase_count[2] ^ phase[245][2]) || (phase_count[3] ^ phase[245][3]) || (phase_count[4] ^ phase[245][4]) || (phase_count[5] ^ phase[245][5]) || (phase_count[6] ^ phase[245][6]) || phase[245][7];
	assign select[246] = (phase_count[0] ^ phase[246][0]) || (phase_count[1] ^ phase[246][1]) || (phase_count[2] ^ phase[246][2]) || (phase_count[3] ^ phase[246][3]) || (phase_count[4] ^ phase[246][4]) || (phase_count[5] ^ phase[246][5]) || (phase_count[6] ^ phase[246][6]) || phase[246][7];
	assign select[247] = (phase_count[0] ^ phase[247][0]) || (phase_count[1] ^ phase[247][1]) || (phase_count[2] ^ phase[247][2]) || (phase_count[3] ^ phase[247][3]) || (phase_count[4] ^ phase[247][4]) || (phase_count[5] ^ phase[247][5]) || (phase_count[6] ^ phase[247][6]) || phase[247][7];
	assign select[248] = (phase_count[0] ^ phase[248][0]) || (phase_count[1] ^ phase[248][1]) || (phase_count[2] ^ phase[248][2]) || (phase_count[3] ^ phase[248][3]) || (phase_count[4] ^ phase[248][4]) || (phase_count[5] ^ phase[248][5]) || (phase_count[6] ^ phase[248][6]) || phase[248][7];
	assign select[249] = (phase_count[0] ^ phase[249][0]) || (phase_count[1] ^ phase[249][1]) || (phase_count[2] ^ phase[249][2]) || (phase_count[3] ^ phase[249][3]) || (phase_count[4] ^ phase[249][4]) || (phase_count[5] ^ phase[249][5]) || (phase_count[6] ^ phase[249][6]) || phase[249][7];
	assign select[250] = (phase_count[0] ^ phase[250][0]) || (phase_count[1] ^ phase[250][1]) || (phase_count[2] ^ phase[250][2]) || (phase_count[3] ^ phase[250][3]) || (phase_count[4] ^ phase[250][4]) || (phase_count[5] ^ phase[250][5]) || (phase_count[6] ^ phase[250][6]) || phase[250][7];
	assign select[251] = (phase_count[0] ^ phase[251][0]) || (phase_count[1] ^ phase[251][1]) || (phase_count[2] ^ phase[251][2]) || (phase_count[3] ^ phase[251][3]) || (phase_count[4] ^ phase[251][4]) || (phase_count[5] ^ phase[251][5]) || (phase_count[6] ^ phase[251][6]) || phase[251][7];
	assign select[252] = (phase_count[0] ^ phase[252][0]) || (phase_count[1] ^ phase[252][1]) || (phase_count[2] ^ phase[252][2]) || (phase_count[3] ^ phase[252][3]) || (phase_count[4] ^ phase[252][4]) || (phase_count[5] ^ phase[252][5]) || (phase_count[6] ^ phase[252][6]) || phase[252][7];
	assign select[253] = (phase_count[0] ^ phase[253][0]) || (phase_count[1] ^ phase[253][1]) || (phase_count[2] ^ phase[253][2]) || (phase_count[3] ^ phase[253][3]) || (phase_count[4] ^ phase[253][4]) || (phase_count[5] ^ phase[253][5]) || (phase_count[6] ^ phase[253][6]) || phase[253][7];
	assign select[254] = (phase_count[0] ^ phase[254][0]) || (phase_count[1] ^ phase[254][1]) || (phase_count[2] ^ phase[254][2]) || (phase_count[3] ^ phase[254][3]) || (phase_count[4] ^ phase[254][4]) || (phase_count[5] ^ phase[254][5]) || (phase_count[6] ^ phase[254][6]) || phase[254][7];
	assign select[255] = (phase_count[0] ^ phase[255][0]) || (phase_count[1] ^ phase[255][1]) || (phase_count[2] ^ phase[255][2]) || (phase_count[3] ^ phase[255][3]) || (phase_count[4] ^ phase[255][4]) || (phase_count[5] ^ phase[255][5]) || (phase_count[6] ^ phase[255][6]) || phase[255][7];
	
	//select_end follows the same logic as select
	//assign select_end[0] = (phase_count[0] ^ phase_end[0][0]) || (phase_count[1] ^ phase_end[0][1]) || (phase_count[2] ^ phase_end[0][2]) || (phase_count[3] ^ phase_end[0][3]) || (phase_count[4] ^ phase_end[0][4]) || (phase_count[5] ^ phase_end[0][5]) || (phase_count[6] ^ phase_end[0][6]) || phase[0][7];
	
	assign select_end[0] = (phase_count[0] ^ phase_end[0][0]) || (phase_count[1] ^ phase_end[0][1]) || (phase_count[2] ^ phase_end[0][2]) || (phase_count[3] ^ phase_end[0][3]) || (phase_count[4] ^ phase_end[0][4]) || (phase_count[5] ^ phase_end[0][5]) || (phase_count[6] ^ phase_end[0][6]) || phase[0][7];
	assign select_end[1] = (phase_count[0] ^ phase_end[1][0]) || (phase_count[1] ^ phase_end[1][1]) || (phase_count[2] ^ phase_end[1][2]) || (phase_count[3] ^ phase_end[1][3]) || (phase_count[4] ^ phase_end[1][4]) || (phase_count[5] ^ phase_end[1][5]) || (phase_count[6] ^ phase_end[1][6]) || phase[1][7];
	assign select_end[2] = (phase_count[0] ^ phase_end[2][0]) || (phase_count[1] ^ phase_end[2][1]) || (phase_count[2] ^ phase_end[2][2]) || (phase_count[3] ^ phase_end[2][3]) || (phase_count[4] ^ phase_end[2][4]) || (phase_count[5] ^ phase_end[2][5]) || (phase_count[6] ^ phase_end[2][6]) || phase[2][7];
	assign select_end[3] = (phase_count[0] ^ phase_end[3][0]) || (phase_count[1] ^ phase_end[3][1]) || (phase_count[2] ^ phase_end[3][2]) || (phase_count[3] ^ phase_end[3][3]) || (phase_count[4] ^ phase_end[3][4]) || (phase_count[5] ^ phase_end[3][5]) || (phase_count[6] ^ phase_end[3][6]) || phase[3][7];
	assign select_end[4] = (phase_count[0] ^ phase_end[4][0]) || (phase_count[1] ^ phase_end[4][1]) || (phase_count[2] ^ phase_end[4][2]) || (phase_count[3] ^ phase_end[4][3]) || (phase_count[4] ^ phase_end[4][4]) || (phase_count[5] ^ phase_end[4][5]) || (phase_count[6] ^ phase_end[4][6]) || phase[4][7];
	assign select_end[5] = (phase_count[0] ^ phase_end[5][0]) || (phase_count[1] ^ phase_end[5][1]) || (phase_count[2] ^ phase_end[5][2]) || (phase_count[3] ^ phase_end[5][3]) || (phase_count[4] ^ phase_end[5][4]) || (phase_count[5] ^ phase_end[5][5]) || (phase_count[6] ^ phase_end[5][6]) || phase[5][7];
	assign select_end[6] = (phase_count[0] ^ phase_end[6][0]) || (phase_count[1] ^ phase_end[6][1]) || (phase_count[2] ^ phase_end[6][2]) || (phase_count[3] ^ phase_end[6][3]) || (phase_count[4] ^ phase_end[6][4]) || (phase_count[5] ^ phase_end[6][5]) || (phase_count[6] ^ phase_end[6][6]) || phase[6][7];
	assign select_end[7] = (phase_count[0] ^ phase_end[7][0]) || (phase_count[1] ^ phase_end[7][1]) || (phase_count[2] ^ phase_end[7][2]) || (phase_count[3] ^ phase_end[7][3]) || (phase_count[4] ^ phase_end[7][4]) || (phase_count[5] ^ phase_end[7][5]) || (phase_count[6] ^ phase_end[7][6]) || phase[7][7];
	assign select_end[8] = (phase_count[0] ^ phase_end[8][0]) || (phase_count[1] ^ phase_end[8][1]) || (phase_count[2] ^ phase_end[8][2]) || (phase_count[3] ^ phase_end[8][3]) || (phase_count[4] ^ phase_end[8][4]) || (phase_count[5] ^ phase_end[8][5]) || (phase_count[6] ^ phase_end[8][6]) || phase[8][7];
	assign select_end[9] = (phase_count[0] ^ phase_end[9][0]) || (phase_count[1] ^ phase_end[9][1]) || (phase_count[2] ^ phase_end[9][2]) || (phase_count[3] ^ phase_end[9][3]) || (phase_count[4] ^ phase_end[9][4]) || (phase_count[5] ^ phase_end[9][5]) || (phase_count[6] ^ phase_end[9][6]) || phase[9][7];
	assign select_end[10] = (phase_count[0] ^ phase_end[10][0]) || (phase_count[1] ^ phase_end[10][1]) || (phase_count[2] ^ phase_end[10][2]) || (phase_count[3] ^ phase_end[10][3]) || (phase_count[4] ^ phase_end[10][4]) || (phase_count[5] ^ phase_end[10][5]) || (phase_count[6] ^ phase_end[10][6]) || phase[10][7];
	assign select_end[11] = (phase_count[0] ^ phase_end[11][0]) || (phase_count[1] ^ phase_end[11][1]) || (phase_count[2] ^ phase_end[11][2]) || (phase_count[3] ^ phase_end[11][3]) || (phase_count[4] ^ phase_end[11][4]) || (phase_count[5] ^ phase_end[11][5]) || (phase_count[6] ^ phase_end[11][6]) || phase[11][7];
	assign select_end[12] = (phase_count[0] ^ phase_end[12][0]) || (phase_count[1] ^ phase_end[12][1]) || (phase_count[2] ^ phase_end[12][2]) || (phase_count[3] ^ phase_end[12][3]) || (phase_count[4] ^ phase_end[12][4]) || (phase_count[5] ^ phase_end[12][5]) || (phase_count[6] ^ phase_end[12][6]) || phase[12][7];
	assign select_end[13] = (phase_count[0] ^ phase_end[13][0]) || (phase_count[1] ^ phase_end[13][1]) || (phase_count[2] ^ phase_end[13][2]) || (phase_count[3] ^ phase_end[13][3]) || (phase_count[4] ^ phase_end[13][4]) || (phase_count[5] ^ phase_end[13][5]) || (phase_count[6] ^ phase_end[13][6]) || phase[13][7];
	assign select_end[14] = (phase_count[0] ^ phase_end[14][0]) || (phase_count[1] ^ phase_end[14][1]) || (phase_count[2] ^ phase_end[14][2]) || (phase_count[3] ^ phase_end[14][3]) || (phase_count[4] ^ phase_end[14][4]) || (phase_count[5] ^ phase_end[14][5]) || (phase_count[6] ^ phase_end[14][6]) || phase[14][7];
	assign select_end[15] = (phase_count[0] ^ phase_end[15][0]) || (phase_count[1] ^ phase_end[15][1]) || (phase_count[2] ^ phase_end[15][2]) || (phase_count[3] ^ phase_end[15][3]) || (phase_count[4] ^ phase_end[15][4]) || (phase_count[5] ^ phase_end[15][5]) || (phase_count[6] ^ phase_end[15][6]) || phase[15][7];
	assign select_end[16] = (phase_count[0] ^ phase_end[16][0]) || (phase_count[1] ^ phase_end[16][1]) || (phase_count[2] ^ phase_end[16][2]) || (phase_count[3] ^ phase_end[16][3]) || (phase_count[4] ^ phase_end[16][4]) || (phase_count[5] ^ phase_end[16][5]) || (phase_count[6] ^ phase_end[16][6]) || phase[16][7];
	assign select_end[17] = (phase_count[0] ^ phase_end[17][0]) || (phase_count[1] ^ phase_end[17][1]) || (phase_count[2] ^ phase_end[17][2]) || (phase_count[3] ^ phase_end[17][3]) || (phase_count[4] ^ phase_end[17][4]) || (phase_count[5] ^ phase_end[17][5]) || (phase_count[6] ^ phase_end[17][6]) || phase[17][7];
	assign select_end[18] = (phase_count[0] ^ phase_end[18][0]) || (phase_count[1] ^ phase_end[18][1]) || (phase_count[2] ^ phase_end[18][2]) || (phase_count[3] ^ phase_end[18][3]) || (phase_count[4] ^ phase_end[18][4]) || (phase_count[5] ^ phase_end[18][5]) || (phase_count[6] ^ phase_end[18][6]) || phase[18][7];
	assign select_end[19] = (phase_count[0] ^ phase_end[19][0]) || (phase_count[1] ^ phase_end[19][1]) || (phase_count[2] ^ phase_end[19][2]) || (phase_count[3] ^ phase_end[19][3]) || (phase_count[4] ^ phase_end[19][4]) || (phase_count[5] ^ phase_end[19][5]) || (phase_count[6] ^ phase_end[19][6]) || phase[19][7];
	assign select_end[20] = (phase_count[0] ^ phase_end[20][0]) || (phase_count[1] ^ phase_end[20][1]) || (phase_count[2] ^ phase_end[20][2]) || (phase_count[3] ^ phase_end[20][3]) || (phase_count[4] ^ phase_end[20][4]) || (phase_count[5] ^ phase_end[20][5]) || (phase_count[6] ^ phase_end[20][6]) || phase[20][7];
	assign select_end[21] = (phase_count[0] ^ phase_end[21][0]) || (phase_count[1] ^ phase_end[21][1]) || (phase_count[2] ^ phase_end[21][2]) || (phase_count[3] ^ phase_end[21][3]) || (phase_count[4] ^ phase_end[21][4]) || (phase_count[5] ^ phase_end[21][5]) || (phase_count[6] ^ phase_end[21][6]) || phase[21][7];
	assign select_end[22] = (phase_count[0] ^ phase_end[22][0]) || (phase_count[1] ^ phase_end[22][1]) || (phase_count[2] ^ phase_end[22][2]) || (phase_count[3] ^ phase_end[22][3]) || (phase_count[4] ^ phase_end[22][4]) || (phase_count[5] ^ phase_end[22][5]) || (phase_count[6] ^ phase_end[22][6]) || phase[22][7];
	assign select_end[23] = (phase_count[0] ^ phase_end[23][0]) || (phase_count[1] ^ phase_end[23][1]) || (phase_count[2] ^ phase_end[23][2]) || (phase_count[3] ^ phase_end[23][3]) || (phase_count[4] ^ phase_end[23][4]) || (phase_count[5] ^ phase_end[23][5]) || (phase_count[6] ^ phase_end[23][6]) || phase[23][7];
	assign select_end[24] = (phase_count[0] ^ phase_end[24][0]) || (phase_count[1] ^ phase_end[24][1]) || (phase_count[2] ^ phase_end[24][2]) || (phase_count[3] ^ phase_end[24][3]) || (phase_count[4] ^ phase_end[24][4]) || (phase_count[5] ^ phase_end[24][5]) || (phase_count[6] ^ phase_end[24][6]) || phase[24][7];
	assign select_end[25] = (phase_count[0] ^ phase_end[25][0]) || (phase_count[1] ^ phase_end[25][1]) || (phase_count[2] ^ phase_end[25][2]) || (phase_count[3] ^ phase_end[25][3]) || (phase_count[4] ^ phase_end[25][4]) || (phase_count[5] ^ phase_end[25][5]) || (phase_count[6] ^ phase_end[25][6]) || phase[25][7];
	assign select_end[26] = (phase_count[0] ^ phase_end[26][0]) || (phase_count[1] ^ phase_end[26][1]) || (phase_count[2] ^ phase_end[26][2]) || (phase_count[3] ^ phase_end[26][3]) || (phase_count[4] ^ phase_end[26][4]) || (phase_count[5] ^ phase_end[26][5]) || (phase_count[6] ^ phase_end[26][6]) || phase[26][7];
	assign select_end[27] = (phase_count[0] ^ phase_end[27][0]) || (phase_count[1] ^ phase_end[27][1]) || (phase_count[2] ^ phase_end[27][2]) || (phase_count[3] ^ phase_end[27][3]) || (phase_count[4] ^ phase_end[27][4]) || (phase_count[5] ^ phase_end[27][5]) || (phase_count[6] ^ phase_end[27][6]) || phase[27][7];
	assign select_end[28] = (phase_count[0] ^ phase_end[28][0]) || (phase_count[1] ^ phase_end[28][1]) || (phase_count[2] ^ phase_end[28][2]) || (phase_count[3] ^ phase_end[28][3]) || (phase_count[4] ^ phase_end[28][4]) || (phase_count[5] ^ phase_end[28][5]) || (phase_count[6] ^ phase_end[28][6]) || phase[28][7];
	assign select_end[29] = (phase_count[0] ^ phase_end[29][0]) || (phase_count[1] ^ phase_end[29][1]) || (phase_count[2] ^ phase_end[29][2]) || (phase_count[3] ^ phase_end[29][3]) || (phase_count[4] ^ phase_end[29][4]) || (phase_count[5] ^ phase_end[29][5]) || (phase_count[6] ^ phase_end[29][6]) || phase[29][7];
	assign select_end[30] = (phase_count[0] ^ phase_end[30][0]) || (phase_count[1] ^ phase_end[30][1]) || (phase_count[2] ^ phase_end[30][2]) || (phase_count[3] ^ phase_end[30][3]) || (phase_count[4] ^ phase_end[30][4]) || (phase_count[5] ^ phase_end[30][5]) || (phase_count[6] ^ phase_end[30][6]) || phase[30][7];
	assign select_end[31] = (phase_count[0] ^ phase_end[31][0]) || (phase_count[1] ^ phase_end[31][1]) || (phase_count[2] ^ phase_end[31][2]) || (phase_count[3] ^ phase_end[31][3]) || (phase_count[4] ^ phase_end[31][4]) || (phase_count[5] ^ phase_end[31][5]) || (phase_count[6] ^ phase_end[31][6]) || phase[31][7];
	assign select_end[32] = (phase_count[0] ^ phase_end[32][0]) || (phase_count[1] ^ phase_end[32][1]) || (phase_count[2] ^ phase_end[32][2]) || (phase_count[3] ^ phase_end[32][3]) || (phase_count[4] ^ phase_end[32][4]) || (phase_count[5] ^ phase_end[32][5]) || (phase_count[6] ^ phase_end[32][6]) || phase[32][7];
	assign select_end[33] = (phase_count[0] ^ phase_end[33][0]) || (phase_count[1] ^ phase_end[33][1]) || (phase_count[2] ^ phase_end[33][2]) || (phase_count[3] ^ phase_end[33][3]) || (phase_count[4] ^ phase_end[33][4]) || (phase_count[5] ^ phase_end[33][5]) || (phase_count[6] ^ phase_end[33][6]) || phase[33][7];
	assign select_end[34] = (phase_count[0] ^ phase_end[34][0]) || (phase_count[1] ^ phase_end[34][1]) || (phase_count[2] ^ phase_end[34][2]) || (phase_count[3] ^ phase_end[34][3]) || (phase_count[4] ^ phase_end[34][4]) || (phase_count[5] ^ phase_end[34][5]) || (phase_count[6] ^ phase_end[34][6]) || phase[34][7];
	assign select_end[35] = (phase_count[0] ^ phase_end[35][0]) || (phase_count[1] ^ phase_end[35][1]) || (phase_count[2] ^ phase_end[35][2]) || (phase_count[3] ^ phase_end[35][3]) || (phase_count[4] ^ phase_end[35][4]) || (phase_count[5] ^ phase_end[35][5]) || (phase_count[6] ^ phase_end[35][6]) || phase[35][7];
	assign select_end[36] = (phase_count[0] ^ phase_end[36][0]) || (phase_count[1] ^ phase_end[36][1]) || (phase_count[2] ^ phase_end[36][2]) || (phase_count[3] ^ phase_end[36][3]) || (phase_count[4] ^ phase_end[36][4]) || (phase_count[5] ^ phase_end[36][5]) || (phase_count[6] ^ phase_end[36][6]) || phase[36][7];
	assign select_end[37] = (phase_count[0] ^ phase_end[37][0]) || (phase_count[1] ^ phase_end[37][1]) || (phase_count[2] ^ phase_end[37][2]) || (phase_count[3] ^ phase_end[37][3]) || (phase_count[4] ^ phase_end[37][4]) || (phase_count[5] ^ phase_end[37][5]) || (phase_count[6] ^ phase_end[37][6]) || phase[37][7];
	assign select_end[38] = (phase_count[0] ^ phase_end[38][0]) || (phase_count[1] ^ phase_end[38][1]) || (phase_count[2] ^ phase_end[38][2]) || (phase_count[3] ^ phase_end[38][3]) || (phase_count[4] ^ phase_end[38][4]) || (phase_count[5] ^ phase_end[38][5]) || (phase_count[6] ^ phase_end[38][6]) || phase[38][7];
	assign select_end[39] = (phase_count[0] ^ phase_end[39][0]) || (phase_count[1] ^ phase_end[39][1]) || (phase_count[2] ^ phase_end[39][2]) || (phase_count[3] ^ phase_end[39][3]) || (phase_count[4] ^ phase_end[39][4]) || (phase_count[5] ^ phase_end[39][5]) || (phase_count[6] ^ phase_end[39][6]) || phase[39][7];
	assign select_end[40] = (phase_count[0] ^ phase_end[40][0]) || (phase_count[1] ^ phase_end[40][1]) || (phase_count[2] ^ phase_end[40][2]) || (phase_count[3] ^ phase_end[40][3]) || (phase_count[4] ^ phase_end[40][4]) || (phase_count[5] ^ phase_end[40][5]) || (phase_count[6] ^ phase_end[40][6]) || phase[40][7];
	assign select_end[41] = (phase_count[0] ^ phase_end[41][0]) || (phase_count[1] ^ phase_end[41][1]) || (phase_count[2] ^ phase_end[41][2]) || (phase_count[3] ^ phase_end[41][3]) || (phase_count[4] ^ phase_end[41][4]) || (phase_count[5] ^ phase_end[41][5]) || (phase_count[6] ^ phase_end[41][6]) || phase[41][7];
	assign select_end[42] = (phase_count[0] ^ phase_end[42][0]) || (phase_count[1] ^ phase_end[42][1]) || (phase_count[2] ^ phase_end[42][2]) || (phase_count[3] ^ phase_end[42][3]) || (phase_count[4] ^ phase_end[42][4]) || (phase_count[5] ^ phase_end[42][5]) || (phase_count[6] ^ phase_end[42][6]) || phase[42][7];
	assign select_end[43] = (phase_count[0] ^ phase_end[43][0]) || (phase_count[1] ^ phase_end[43][1]) || (phase_count[2] ^ phase_end[43][2]) || (phase_count[3] ^ phase_end[43][3]) || (phase_count[4] ^ phase_end[43][4]) || (phase_count[5] ^ phase_end[43][5]) || (phase_count[6] ^ phase_end[43][6]) || phase[43][7];
	assign select_end[44] = (phase_count[0] ^ phase_end[44][0]) || (phase_count[1] ^ phase_end[44][1]) || (phase_count[2] ^ phase_end[44][2]) || (phase_count[3] ^ phase_end[44][3]) || (phase_count[4] ^ phase_end[44][4]) || (phase_count[5] ^ phase_end[44][5]) || (phase_count[6] ^ phase_end[44][6]) || phase[44][7];
	assign select_end[45] = (phase_count[0] ^ phase_end[45][0]) || (phase_count[1] ^ phase_end[45][1]) || (phase_count[2] ^ phase_end[45][2]) || (phase_count[3] ^ phase_end[45][3]) || (phase_count[4] ^ phase_end[45][4]) || (phase_count[5] ^ phase_end[45][5]) || (phase_count[6] ^ phase_end[45][6]) || phase[45][7];
	assign select_end[46] = (phase_count[0] ^ phase_end[46][0]) || (phase_count[1] ^ phase_end[46][1]) || (phase_count[2] ^ phase_end[46][2]) || (phase_count[3] ^ phase_end[46][3]) || (phase_count[4] ^ phase_end[46][4]) || (phase_count[5] ^ phase_end[46][5]) || (phase_count[6] ^ phase_end[46][6]) || phase[46][7];
	assign select_end[47] = (phase_count[0] ^ phase_end[47][0]) || (phase_count[1] ^ phase_end[47][1]) || (phase_count[2] ^ phase_end[47][2]) || (phase_count[3] ^ phase_end[47][3]) || (phase_count[4] ^ phase_end[47][4]) || (phase_count[5] ^ phase_end[47][5]) || (phase_count[6] ^ phase_end[47][6]) || phase[47][7];
	assign select_end[48] = (phase_count[0] ^ phase_end[48][0]) || (phase_count[1] ^ phase_end[48][1]) || (phase_count[2] ^ phase_end[48][2]) || (phase_count[3] ^ phase_end[48][3]) || (phase_count[4] ^ phase_end[48][4]) || (phase_count[5] ^ phase_end[48][5]) || (phase_count[6] ^ phase_end[48][6]) || phase[48][7];
	assign select_end[49] = (phase_count[0] ^ phase_end[49][0]) || (phase_count[1] ^ phase_end[49][1]) || (phase_count[2] ^ phase_end[49][2]) || (phase_count[3] ^ phase_end[49][3]) || (phase_count[4] ^ phase_end[49][4]) || (phase_count[5] ^ phase_end[49][5]) || (phase_count[6] ^ phase_end[49][6]) || phase[49][7];
	assign select_end[50] = (phase_count[0] ^ phase_end[50][0]) || (phase_count[1] ^ phase_end[50][1]) || (phase_count[2] ^ phase_end[50][2]) || (phase_count[3] ^ phase_end[50][3]) || (phase_count[4] ^ phase_end[50][4]) || (phase_count[5] ^ phase_end[50][5]) || (phase_count[6] ^ phase_end[50][6]) || phase[50][7];
	assign select_end[51] = (phase_count[0] ^ phase_end[51][0]) || (phase_count[1] ^ phase_end[51][1]) || (phase_count[2] ^ phase_end[51][2]) || (phase_count[3] ^ phase_end[51][3]) || (phase_count[4] ^ phase_end[51][4]) || (phase_count[5] ^ phase_end[51][5]) || (phase_count[6] ^ phase_end[51][6]) || phase[51][7];
	assign select_end[52] = (phase_count[0] ^ phase_end[52][0]) || (phase_count[1] ^ phase_end[52][1]) || (phase_count[2] ^ phase_end[52][2]) || (phase_count[3] ^ phase_end[52][3]) || (phase_count[4] ^ phase_end[52][4]) || (phase_count[5] ^ phase_end[52][5]) || (phase_count[6] ^ phase_end[52][6]) || phase[52][7];
	assign select_end[53] = (phase_count[0] ^ phase_end[53][0]) || (phase_count[1] ^ phase_end[53][1]) || (phase_count[2] ^ phase_end[53][2]) || (phase_count[3] ^ phase_end[53][3]) || (phase_count[4] ^ phase_end[53][4]) || (phase_count[5] ^ phase_end[53][5]) || (phase_count[6] ^ phase_end[53][6]) || phase[53][7];
	assign select_end[54] = (phase_count[0] ^ phase_end[54][0]) || (phase_count[1] ^ phase_end[54][1]) || (phase_count[2] ^ phase_end[54][2]) || (phase_count[3] ^ phase_end[54][3]) || (phase_count[4] ^ phase_end[54][4]) || (phase_count[5] ^ phase_end[54][5]) || (phase_count[6] ^ phase_end[54][6]) || phase[54][7];
	assign select_end[55] = (phase_count[0] ^ phase_end[55][0]) || (phase_count[1] ^ phase_end[55][1]) || (phase_count[2] ^ phase_end[55][2]) || (phase_count[3] ^ phase_end[55][3]) || (phase_count[4] ^ phase_end[55][4]) || (phase_count[5] ^ phase_end[55][5]) || (phase_count[6] ^ phase_end[55][6]) || phase[55][7];
	assign select_end[56] = (phase_count[0] ^ phase_end[56][0]) || (phase_count[1] ^ phase_end[56][1]) || (phase_count[2] ^ phase_end[56][2]) || (phase_count[3] ^ phase_end[56][3]) || (phase_count[4] ^ phase_end[56][4]) || (phase_count[5] ^ phase_end[56][5]) || (phase_count[6] ^ phase_end[56][6]) || phase[56][7];
	assign select_end[57] = (phase_count[0] ^ phase_end[57][0]) || (phase_count[1] ^ phase_end[57][1]) || (phase_count[2] ^ phase_end[57][2]) || (phase_count[3] ^ phase_end[57][3]) || (phase_count[4] ^ phase_end[57][4]) || (phase_count[5] ^ phase_end[57][5]) || (phase_count[6] ^ phase_end[57][6]) || phase[57][7];
	assign select_end[58] = (phase_count[0] ^ phase_end[58][0]) || (phase_count[1] ^ phase_end[58][1]) || (phase_count[2] ^ phase_end[58][2]) || (phase_count[3] ^ phase_end[58][3]) || (phase_count[4] ^ phase_end[58][4]) || (phase_count[5] ^ phase_end[58][5]) || (phase_count[6] ^ phase_end[58][6]) || phase[58][7];
	assign select_end[59] = (phase_count[0] ^ phase_end[59][0]) || (phase_count[1] ^ phase_end[59][1]) || (phase_count[2] ^ phase_end[59][2]) || (phase_count[3] ^ phase_end[59][3]) || (phase_count[4] ^ phase_end[59][4]) || (phase_count[5] ^ phase_end[59][5]) || (phase_count[6] ^ phase_end[59][6]) || phase[59][7];
	assign select_end[60] = (phase_count[0] ^ phase_end[60][0]) || (phase_count[1] ^ phase_end[60][1]) || (phase_count[2] ^ phase_end[60][2]) || (phase_count[3] ^ phase_end[60][3]) || (phase_count[4] ^ phase_end[60][4]) || (phase_count[5] ^ phase_end[60][5]) || (phase_count[6] ^ phase_end[60][6]) || phase[60][7];
	assign select_end[61] = (phase_count[0] ^ phase_end[61][0]) || (phase_count[1] ^ phase_end[61][1]) || (phase_count[2] ^ phase_end[61][2]) || (phase_count[3] ^ phase_end[61][3]) || (phase_count[4] ^ phase_end[61][4]) || (phase_count[5] ^ phase_end[61][5]) || (phase_count[6] ^ phase_end[61][6]) || phase[61][7];
	assign select_end[62] = (phase_count[0] ^ phase_end[62][0]) || (phase_count[1] ^ phase_end[62][1]) || (phase_count[2] ^ phase_end[62][2]) || (phase_count[3] ^ phase_end[62][3]) || (phase_count[4] ^ phase_end[62][4]) || (phase_count[5] ^ phase_end[62][5]) || (phase_count[6] ^ phase_end[62][6]) || phase[62][7];
	assign select_end[63] = (phase_count[0] ^ phase_end[63][0]) || (phase_count[1] ^ phase_end[63][1]) || (phase_count[2] ^ phase_end[63][2]) || (phase_count[3] ^ phase_end[63][3]) || (phase_count[4] ^ phase_end[63][4]) || (phase_count[5] ^ phase_end[63][5]) || (phase_count[6] ^ phase_end[63][6]) || phase[63][7];
	assign select_end[64] = (phase_count[0] ^ phase_end[64][0]) || (phase_count[1] ^ phase_end[64][1]) || (phase_count[2] ^ phase_end[64][2]) || (phase_count[3] ^ phase_end[64][3]) || (phase_count[4] ^ phase_end[64][4]) || (phase_count[5] ^ phase_end[64][5]) || (phase_count[6] ^ phase_end[64][6]) || phase[64][7];
	assign select_end[65] = (phase_count[0] ^ phase_end[65][0]) || (phase_count[1] ^ phase_end[65][1]) || (phase_count[2] ^ phase_end[65][2]) || (phase_count[3] ^ phase_end[65][3]) || (phase_count[4] ^ phase_end[65][4]) || (phase_count[5] ^ phase_end[65][5]) || (phase_count[6] ^ phase_end[65][6]) || phase[65][7];
	assign select_end[66] = (phase_count[0] ^ phase_end[66][0]) || (phase_count[1] ^ phase_end[66][1]) || (phase_count[2] ^ phase_end[66][2]) || (phase_count[3] ^ phase_end[66][3]) || (phase_count[4] ^ phase_end[66][4]) || (phase_count[5] ^ phase_end[66][5]) || (phase_count[6] ^ phase_end[66][6]) || phase[66][7];
	assign select_end[67] = (phase_count[0] ^ phase_end[67][0]) || (phase_count[1] ^ phase_end[67][1]) || (phase_count[2] ^ phase_end[67][2]) || (phase_count[3] ^ phase_end[67][3]) || (phase_count[4] ^ phase_end[67][4]) || (phase_count[5] ^ phase_end[67][5]) || (phase_count[6] ^ phase_end[67][6]) || phase[67][7];
	assign select_end[68] = (phase_count[0] ^ phase_end[68][0]) || (phase_count[1] ^ phase_end[68][1]) || (phase_count[2] ^ phase_end[68][2]) || (phase_count[3] ^ phase_end[68][3]) || (phase_count[4] ^ phase_end[68][4]) || (phase_count[5] ^ phase_end[68][5]) || (phase_count[6] ^ phase_end[68][6]) || phase[68][7];
	assign select_end[69] = (phase_count[0] ^ phase_end[69][0]) || (phase_count[1] ^ phase_end[69][1]) || (phase_count[2] ^ phase_end[69][2]) || (phase_count[3] ^ phase_end[69][3]) || (phase_count[4] ^ phase_end[69][4]) || (phase_count[5] ^ phase_end[69][5]) || (phase_count[6] ^ phase_end[69][6]) || phase[69][7];
	assign select_end[70] = (phase_count[0] ^ phase_end[70][0]) || (phase_count[1] ^ phase_end[70][1]) || (phase_count[2] ^ phase_end[70][2]) || (phase_count[3] ^ phase_end[70][3]) || (phase_count[4] ^ phase_end[70][4]) || (phase_count[5] ^ phase_end[70][5]) || (phase_count[6] ^ phase_end[70][6]) || phase[70][7];
	assign select_end[71] = (phase_count[0] ^ phase_end[71][0]) || (phase_count[1] ^ phase_end[71][1]) || (phase_count[2] ^ phase_end[71][2]) || (phase_count[3] ^ phase_end[71][3]) || (phase_count[4] ^ phase_end[71][4]) || (phase_count[5] ^ phase_end[71][5]) || (phase_count[6] ^ phase_end[71][6]) || phase[71][7];
	assign select_end[72] = (phase_count[0] ^ phase_end[72][0]) || (phase_count[1] ^ phase_end[72][1]) || (phase_count[2] ^ phase_end[72][2]) || (phase_count[3] ^ phase_end[72][3]) || (phase_count[4] ^ phase_end[72][4]) || (phase_count[5] ^ phase_end[72][5]) || (phase_count[6] ^ phase_end[72][6]) || phase[72][7];
	assign select_end[73] = (phase_count[0] ^ phase_end[73][0]) || (phase_count[1] ^ phase_end[73][1]) || (phase_count[2] ^ phase_end[73][2]) || (phase_count[3] ^ phase_end[73][3]) || (phase_count[4] ^ phase_end[73][4]) || (phase_count[5] ^ phase_end[73][5]) || (phase_count[6] ^ phase_end[73][6]) || phase[73][7];
	assign select_end[74] = (phase_count[0] ^ phase_end[74][0]) || (phase_count[1] ^ phase_end[74][1]) || (phase_count[2] ^ phase_end[74][2]) || (phase_count[3] ^ phase_end[74][3]) || (phase_count[4] ^ phase_end[74][4]) || (phase_count[5] ^ phase_end[74][5]) || (phase_count[6] ^ phase_end[74][6]) || phase[74][7];
	assign select_end[75] = (phase_count[0] ^ phase_end[75][0]) || (phase_count[1] ^ phase_end[75][1]) || (phase_count[2] ^ phase_end[75][2]) || (phase_count[3] ^ phase_end[75][3]) || (phase_count[4] ^ phase_end[75][4]) || (phase_count[5] ^ phase_end[75][5]) || (phase_count[6] ^ phase_end[75][6]) || phase[75][7];
	assign select_end[76] = (phase_count[0] ^ phase_end[76][0]) || (phase_count[1] ^ phase_end[76][1]) || (phase_count[2] ^ phase_end[76][2]) || (phase_count[3] ^ phase_end[76][3]) || (phase_count[4] ^ phase_end[76][4]) || (phase_count[5] ^ phase_end[76][5]) || (phase_count[6] ^ phase_end[76][6]) || phase[76][7];
	assign select_end[77] = (phase_count[0] ^ phase_end[77][0]) || (phase_count[1] ^ phase_end[77][1]) || (phase_count[2] ^ phase_end[77][2]) || (phase_count[3] ^ phase_end[77][3]) || (phase_count[4] ^ phase_end[77][4]) || (phase_count[5] ^ phase_end[77][5]) || (phase_count[6] ^ phase_end[77][6]) || phase[77][7];
	assign select_end[78] = (phase_count[0] ^ phase_end[78][0]) || (phase_count[1] ^ phase_end[78][1]) || (phase_count[2] ^ phase_end[78][2]) || (phase_count[3] ^ phase_end[78][3]) || (phase_count[4] ^ phase_end[78][4]) || (phase_count[5] ^ phase_end[78][5]) || (phase_count[6] ^ phase_end[78][6]) || phase[78][7];
	assign select_end[79] = (phase_count[0] ^ phase_end[79][0]) || (phase_count[1] ^ phase_end[79][1]) || (phase_count[2] ^ phase_end[79][2]) || (phase_count[3] ^ phase_end[79][3]) || (phase_count[4] ^ phase_end[79][4]) || (phase_count[5] ^ phase_end[79][5]) || (phase_count[6] ^ phase_end[79][6]) || phase[79][7];
	assign select_end[80] = (phase_count[0] ^ phase_end[80][0]) || (phase_count[1] ^ phase_end[80][1]) || (phase_count[2] ^ phase_end[80][2]) || (phase_count[3] ^ phase_end[80][3]) || (phase_count[4] ^ phase_end[80][4]) || (phase_count[5] ^ phase_end[80][5]) || (phase_count[6] ^ phase_end[80][6]) || phase[80][7];
	assign select_end[81] = (phase_count[0] ^ phase_end[81][0]) || (phase_count[1] ^ phase_end[81][1]) || (phase_count[2] ^ phase_end[81][2]) || (phase_count[3] ^ phase_end[81][3]) || (phase_count[4] ^ phase_end[81][4]) || (phase_count[5] ^ phase_end[81][5]) || (phase_count[6] ^ phase_end[81][6]) || phase[81][7];
	assign select_end[82] = (phase_count[0] ^ phase_end[82][0]) || (phase_count[1] ^ phase_end[82][1]) || (phase_count[2] ^ phase_end[82][2]) || (phase_count[3] ^ phase_end[82][3]) || (phase_count[4] ^ phase_end[82][4]) || (phase_count[5] ^ phase_end[82][5]) || (phase_count[6] ^ phase_end[82][6]) || phase[82][7];
	assign select_end[83] = (phase_count[0] ^ phase_end[83][0]) || (phase_count[1] ^ phase_end[83][1]) || (phase_count[2] ^ phase_end[83][2]) || (phase_count[3] ^ phase_end[83][3]) || (phase_count[4] ^ phase_end[83][4]) || (phase_count[5] ^ phase_end[83][5]) || (phase_count[6] ^ phase_end[83][6]) || phase[83][7];
	assign select_end[84] = (phase_count[0] ^ phase_end[84][0]) || (phase_count[1] ^ phase_end[84][1]) || (phase_count[2] ^ phase_end[84][2]) || (phase_count[3] ^ phase_end[84][3]) || (phase_count[4] ^ phase_end[84][4]) || (phase_count[5] ^ phase_end[84][5]) || (phase_count[6] ^ phase_end[84][6]) || phase[84][7];
	assign select_end[85] = (phase_count[0] ^ phase_end[85][0]) || (phase_count[1] ^ phase_end[85][1]) || (phase_count[2] ^ phase_end[85][2]) || (phase_count[3] ^ phase_end[85][3]) || (phase_count[4] ^ phase_end[85][4]) || (phase_count[5] ^ phase_end[85][5]) || (phase_count[6] ^ phase_end[85][6]) || phase[85][7];
	assign select_end[86] = (phase_count[0] ^ phase_end[86][0]) || (phase_count[1] ^ phase_end[86][1]) || (phase_count[2] ^ phase_end[86][2]) || (phase_count[3] ^ phase_end[86][3]) || (phase_count[4] ^ phase_end[86][4]) || (phase_count[5] ^ phase_end[86][5]) || (phase_count[6] ^ phase_end[86][6]) || phase[86][7];
	assign select_end[87] = (phase_count[0] ^ phase_end[87][0]) || (phase_count[1] ^ phase_end[87][1]) || (phase_count[2] ^ phase_end[87][2]) || (phase_count[3] ^ phase_end[87][3]) || (phase_count[4] ^ phase_end[87][4]) || (phase_count[5] ^ phase_end[87][5]) || (phase_count[6] ^ phase_end[87][6]) || phase[87][7];
	assign select_end[88] = (phase_count[0] ^ phase_end[88][0]) || (phase_count[1] ^ phase_end[88][1]) || (phase_count[2] ^ phase_end[88][2]) || (phase_count[3] ^ phase_end[88][3]) || (phase_count[4] ^ phase_end[88][4]) || (phase_count[5] ^ phase_end[88][5]) || (phase_count[6] ^ phase_end[88][6]) || phase[88][7];
	assign select_end[89] = (phase_count[0] ^ phase_end[89][0]) || (phase_count[1] ^ phase_end[89][1]) || (phase_count[2] ^ phase_end[89][2]) || (phase_count[3] ^ phase_end[89][3]) || (phase_count[4] ^ phase_end[89][4]) || (phase_count[5] ^ phase_end[89][5]) || (phase_count[6] ^ phase_end[89][6]) || phase[89][7];
	assign select_end[90] = (phase_count[0] ^ phase_end[90][0]) || (phase_count[1] ^ phase_end[90][1]) || (phase_count[2] ^ phase_end[90][2]) || (phase_count[3] ^ phase_end[90][3]) || (phase_count[4] ^ phase_end[90][4]) || (phase_count[5] ^ phase_end[90][5]) || (phase_count[6] ^ phase_end[90][6]) || phase[90][7];
	assign select_end[91] = (phase_count[0] ^ phase_end[91][0]) || (phase_count[1] ^ phase_end[91][1]) || (phase_count[2] ^ phase_end[91][2]) || (phase_count[3] ^ phase_end[91][3]) || (phase_count[4] ^ phase_end[91][4]) || (phase_count[5] ^ phase_end[91][5]) || (phase_count[6] ^ phase_end[91][6]) || phase[91][7];
	assign select_end[92] = (phase_count[0] ^ phase_end[92][0]) || (phase_count[1] ^ phase_end[92][1]) || (phase_count[2] ^ phase_end[92][2]) || (phase_count[3] ^ phase_end[92][3]) || (phase_count[4] ^ phase_end[92][4]) || (phase_count[5] ^ phase_end[92][5]) || (phase_count[6] ^ phase_end[92][6]) || phase[92][7];
	assign select_end[93] = (phase_count[0] ^ phase_end[93][0]) || (phase_count[1] ^ phase_end[93][1]) || (phase_count[2] ^ phase_end[93][2]) || (phase_count[3] ^ phase_end[93][3]) || (phase_count[4] ^ phase_end[93][4]) || (phase_count[5] ^ phase_end[93][5]) || (phase_count[6] ^ phase_end[93][6]) || phase[93][7];
	assign select_end[94] = (phase_count[0] ^ phase_end[94][0]) || (phase_count[1] ^ phase_end[94][1]) || (phase_count[2] ^ phase_end[94][2]) || (phase_count[3] ^ phase_end[94][3]) || (phase_count[4] ^ phase_end[94][4]) || (phase_count[5] ^ phase_end[94][5]) || (phase_count[6] ^ phase_end[94][6]) || phase[94][7];
	assign select_end[95] = (phase_count[0] ^ phase_end[95][0]) || (phase_count[1] ^ phase_end[95][1]) || (phase_count[2] ^ phase_end[95][2]) || (phase_count[3] ^ phase_end[95][3]) || (phase_count[4] ^ phase_end[95][4]) || (phase_count[5] ^ phase_end[95][5]) || (phase_count[6] ^ phase_end[95][6]) || phase[95][7];
	assign select_end[96] = (phase_count[0] ^ phase_end[96][0]) || (phase_count[1] ^ phase_end[96][1]) || (phase_count[2] ^ phase_end[96][2]) || (phase_count[3] ^ phase_end[96][3]) || (phase_count[4] ^ phase_end[96][4]) || (phase_count[5] ^ phase_end[96][5]) || (phase_count[6] ^ phase_end[96][6]) || phase[96][7];
	assign select_end[97] = (phase_count[0] ^ phase_end[97][0]) || (phase_count[1] ^ phase_end[97][1]) || (phase_count[2] ^ phase_end[97][2]) || (phase_count[3] ^ phase_end[97][3]) || (phase_count[4] ^ phase_end[97][4]) || (phase_count[5] ^ phase_end[97][5]) || (phase_count[6] ^ phase_end[97][6]) || phase[97][7];
	assign select_end[98] = (phase_count[0] ^ phase_end[98][0]) || (phase_count[1] ^ phase_end[98][1]) || (phase_count[2] ^ phase_end[98][2]) || (phase_count[3] ^ phase_end[98][3]) || (phase_count[4] ^ phase_end[98][4]) || (phase_count[5] ^ phase_end[98][5]) || (phase_count[6] ^ phase_end[98][6]) || phase[98][7];
	assign select_end[99] = (phase_count[0] ^ phase_end[99][0]) || (phase_count[1] ^ phase_end[99][1]) || (phase_count[2] ^ phase_end[99][2]) || (phase_count[3] ^ phase_end[99][3]) || (phase_count[4] ^ phase_end[99][4]) || (phase_count[5] ^ phase_end[99][5]) || (phase_count[6] ^ phase_end[99][6]) || phase[99][7];
	assign select_end[100] = (phase_count[0] ^ phase_end[100][0]) || (phase_count[1] ^ phase_end[100][1]) || (phase_count[2] ^ phase_end[100][2]) || (phase_count[3] ^ phase_end[100][3]) || (phase_count[4] ^ phase_end[100][4]) || (phase_count[5] ^ phase_end[100][5]) || (phase_count[6] ^ phase_end[100][6]) || phase[100][7];
	assign select_end[101] = (phase_count[0] ^ phase_end[101][0]) || (phase_count[1] ^ phase_end[101][1]) || (phase_count[2] ^ phase_end[101][2]) || (phase_count[3] ^ phase_end[101][3]) || (phase_count[4] ^ phase_end[101][4]) || (phase_count[5] ^ phase_end[101][5]) || (phase_count[6] ^ phase_end[101][6]) || phase[101][7];
	assign select_end[102] = (phase_count[0] ^ phase_end[102][0]) || (phase_count[1] ^ phase_end[102][1]) || (phase_count[2] ^ phase_end[102][2]) || (phase_count[3] ^ phase_end[102][3]) || (phase_count[4] ^ phase_end[102][4]) || (phase_count[5] ^ phase_end[102][5]) || (phase_count[6] ^ phase_end[102][6]) || phase[102][7];
	assign select_end[103] = (phase_count[0] ^ phase_end[103][0]) || (phase_count[1] ^ phase_end[103][1]) || (phase_count[2] ^ phase_end[103][2]) || (phase_count[3] ^ phase_end[103][3]) || (phase_count[4] ^ phase_end[103][4]) || (phase_count[5] ^ phase_end[103][5]) || (phase_count[6] ^ phase_end[103][6]) || phase[103][7];
	assign select_end[104] = (phase_count[0] ^ phase_end[104][0]) || (phase_count[1] ^ phase_end[104][1]) || (phase_count[2] ^ phase_end[104][2]) || (phase_count[3] ^ phase_end[104][3]) || (phase_count[4] ^ phase_end[104][4]) || (phase_count[5] ^ phase_end[104][5]) || (phase_count[6] ^ phase_end[104][6]) || phase[104][7];
	assign select_end[105] = (phase_count[0] ^ phase_end[105][0]) || (phase_count[1] ^ phase_end[105][1]) || (phase_count[2] ^ phase_end[105][2]) || (phase_count[3] ^ phase_end[105][3]) || (phase_count[4] ^ phase_end[105][4]) || (phase_count[5] ^ phase_end[105][5]) || (phase_count[6] ^ phase_end[105][6]) || phase[105][7];
	assign select_end[106] = (phase_count[0] ^ phase_end[106][0]) || (phase_count[1] ^ phase_end[106][1]) || (phase_count[2] ^ phase_end[106][2]) || (phase_count[3] ^ phase_end[106][3]) || (phase_count[4] ^ phase_end[106][4]) || (phase_count[5] ^ phase_end[106][5]) || (phase_count[6] ^ phase_end[106][6]) || phase[106][7];
	assign select_end[107] = (phase_count[0] ^ phase_end[107][0]) || (phase_count[1] ^ phase_end[107][1]) || (phase_count[2] ^ phase_end[107][2]) || (phase_count[3] ^ phase_end[107][3]) || (phase_count[4] ^ phase_end[107][4]) || (phase_count[5] ^ phase_end[107][5]) || (phase_count[6] ^ phase_end[107][6]) || phase[107][7];
	assign select_end[108] = (phase_count[0] ^ phase_end[108][0]) || (phase_count[1] ^ phase_end[108][1]) || (phase_count[2] ^ phase_end[108][2]) || (phase_count[3] ^ phase_end[108][3]) || (phase_count[4] ^ phase_end[108][4]) || (phase_count[5] ^ phase_end[108][5]) || (phase_count[6] ^ phase_end[108][6]) || phase[108][7];
	assign select_end[109] = (phase_count[0] ^ phase_end[109][0]) || (phase_count[1] ^ phase_end[109][1]) || (phase_count[2] ^ phase_end[109][2]) || (phase_count[3] ^ phase_end[109][3]) || (phase_count[4] ^ phase_end[109][4]) || (phase_count[5] ^ phase_end[109][5]) || (phase_count[6] ^ phase_end[109][6]) || phase[109][7];
	assign select_end[110] = (phase_count[0] ^ phase_end[110][0]) || (phase_count[1] ^ phase_end[110][1]) || (phase_count[2] ^ phase_end[110][2]) || (phase_count[3] ^ phase_end[110][3]) || (phase_count[4] ^ phase_end[110][4]) || (phase_count[5] ^ phase_end[110][5]) || (phase_count[6] ^ phase_end[110][6]) || phase[110][7];
	assign select_end[111] = (phase_count[0] ^ phase_end[111][0]) || (phase_count[1] ^ phase_end[111][1]) || (phase_count[2] ^ phase_end[111][2]) || (phase_count[3] ^ phase_end[111][3]) || (phase_count[4] ^ phase_end[111][4]) || (phase_count[5] ^ phase_end[111][5]) || (phase_count[6] ^ phase_end[111][6]) || phase[111][7];
	assign select_end[112] = (phase_count[0] ^ phase_end[112][0]) || (phase_count[1] ^ phase_end[112][1]) || (phase_count[2] ^ phase_end[112][2]) || (phase_count[3] ^ phase_end[112][3]) || (phase_count[4] ^ phase_end[112][4]) || (phase_count[5] ^ phase_end[112][5]) || (phase_count[6] ^ phase_end[112][6]) || phase[112][7];
	assign select_end[113] = (phase_count[0] ^ phase_end[113][0]) || (phase_count[1] ^ phase_end[113][1]) || (phase_count[2] ^ phase_end[113][2]) || (phase_count[3] ^ phase_end[113][3]) || (phase_count[4] ^ phase_end[113][4]) || (phase_count[5] ^ phase_end[113][5]) || (phase_count[6] ^ phase_end[113][6]) || phase[113][7];
	assign select_end[114] = (phase_count[0] ^ phase_end[114][0]) || (phase_count[1] ^ phase_end[114][1]) || (phase_count[2] ^ phase_end[114][2]) || (phase_count[3] ^ phase_end[114][3]) || (phase_count[4] ^ phase_end[114][4]) || (phase_count[5] ^ phase_end[114][5]) || (phase_count[6] ^ phase_end[114][6]) || phase[114][7];
	assign select_end[115] = (phase_count[0] ^ phase_end[115][0]) || (phase_count[1] ^ phase_end[115][1]) || (phase_count[2] ^ phase_end[115][2]) || (phase_count[3] ^ phase_end[115][3]) || (phase_count[4] ^ phase_end[115][4]) || (phase_count[5] ^ phase_end[115][5]) || (phase_count[6] ^ phase_end[115][6]) || phase[115][7];
	assign select_end[116] = (phase_count[0] ^ phase_end[116][0]) || (phase_count[1] ^ phase_end[116][1]) || (phase_count[2] ^ phase_end[116][2]) || (phase_count[3] ^ phase_end[116][3]) || (phase_count[4] ^ phase_end[116][4]) || (phase_count[5] ^ phase_end[116][5]) || (phase_count[6] ^ phase_end[116][6]) || phase[116][7];
	assign select_end[117] = (phase_count[0] ^ phase_end[117][0]) || (phase_count[1] ^ phase_end[117][1]) || (phase_count[2] ^ phase_end[117][2]) || (phase_count[3] ^ phase_end[117][3]) || (phase_count[4] ^ phase_end[117][4]) || (phase_count[5] ^ phase_end[117][5]) || (phase_count[6] ^ phase_end[117][6]) || phase[117][7];
	assign select_end[118] = (phase_count[0] ^ phase_end[118][0]) || (phase_count[1] ^ phase_end[118][1]) || (phase_count[2] ^ phase_end[118][2]) || (phase_count[3] ^ phase_end[118][3]) || (phase_count[4] ^ phase_end[118][4]) || (phase_count[5] ^ phase_end[118][5]) || (phase_count[6] ^ phase_end[118][6]) || phase[118][7];
	assign select_end[119] = (phase_count[0] ^ phase_end[119][0]) || (phase_count[1] ^ phase_end[119][1]) || (phase_count[2] ^ phase_end[119][2]) || (phase_count[3] ^ phase_end[119][3]) || (phase_count[4] ^ phase_end[119][4]) || (phase_count[5] ^ phase_end[119][5]) || (phase_count[6] ^ phase_end[119][6]) || phase[119][7];
	assign select_end[120] = (phase_count[0] ^ phase_end[120][0]) || (phase_count[1] ^ phase_end[120][1]) || (phase_count[2] ^ phase_end[120][2]) || (phase_count[3] ^ phase_end[120][3]) || (phase_count[4] ^ phase_end[120][4]) || (phase_count[5] ^ phase_end[120][5]) || (phase_count[6] ^ phase_end[120][6]) || phase[120][7];
	assign select_end[121] = (phase_count[0] ^ phase_end[121][0]) || (phase_count[1] ^ phase_end[121][1]) || (phase_count[2] ^ phase_end[121][2]) || (phase_count[3] ^ phase_end[121][3]) || (phase_count[4] ^ phase_end[121][4]) || (phase_count[5] ^ phase_end[121][5]) || (phase_count[6] ^ phase_end[121][6]) || phase[121][7];
	assign select_end[122] = (phase_count[0] ^ phase_end[122][0]) || (phase_count[1] ^ phase_end[122][1]) || (phase_count[2] ^ phase_end[122][2]) || (phase_count[3] ^ phase_end[122][3]) || (phase_count[4] ^ phase_end[122][4]) || (phase_count[5] ^ phase_end[122][5]) || (phase_count[6] ^ phase_end[122][6]) || phase[122][7];
	assign select_end[123] = (phase_count[0] ^ phase_end[123][0]) || (phase_count[1] ^ phase_end[123][1]) || (phase_count[2] ^ phase_end[123][2]) || (phase_count[3] ^ phase_end[123][3]) || (phase_count[4] ^ phase_end[123][4]) || (phase_count[5] ^ phase_end[123][5]) || (phase_count[6] ^ phase_end[123][6]) || phase[123][7];
	assign select_end[124] = (phase_count[0] ^ phase_end[124][0]) || (phase_count[1] ^ phase_end[124][1]) || (phase_count[2] ^ phase_end[124][2]) || (phase_count[3] ^ phase_end[124][3]) || (phase_count[4] ^ phase_end[124][4]) || (phase_count[5] ^ phase_end[124][5]) || (phase_count[6] ^ phase_end[124][6]) || phase[124][7];
	assign select_end[125] = (phase_count[0] ^ phase_end[125][0]) || (phase_count[1] ^ phase_end[125][1]) || (phase_count[2] ^ phase_end[125][2]) || (phase_count[3] ^ phase_end[125][3]) || (phase_count[4] ^ phase_end[125][4]) || (phase_count[5] ^ phase_end[125][5]) || (phase_count[6] ^ phase_end[125][6]) || phase[125][7];
	assign select_end[126] = (phase_count[0] ^ phase_end[126][0]) || (phase_count[1] ^ phase_end[126][1]) || (phase_count[2] ^ phase_end[126][2]) || (phase_count[3] ^ phase_end[126][3]) || (phase_count[4] ^ phase_end[126][4]) || (phase_count[5] ^ phase_end[126][5]) || (phase_count[6] ^ phase_end[126][6]) || phase[126][7];
	assign select_end[127] = (phase_count[0] ^ phase_end[127][0]) || (phase_count[1] ^ phase_end[127][1]) || (phase_count[2] ^ phase_end[127][2]) || (phase_count[3] ^ phase_end[127][3]) || (phase_count[4] ^ phase_end[127][4]) || (phase_count[5] ^ phase_end[127][5]) || (phase_count[6] ^ phase_end[127][6]) || phase[127][7];
	assign select_end[128] = (phase_count[0] ^ phase_end[128][0]) || (phase_count[1] ^ phase_end[128][1]) || (phase_count[2] ^ phase_end[128][2]) || (phase_count[3] ^ phase_end[128][3]) || (phase_count[4] ^ phase_end[128][4]) || (phase_count[5] ^ phase_end[128][5]) || (phase_count[6] ^ phase_end[128][6]) || phase[128][7];
	assign select_end[129] = (phase_count[0] ^ phase_end[129][0]) || (phase_count[1] ^ phase_end[129][1]) || (phase_count[2] ^ phase_end[129][2]) || (phase_count[3] ^ phase_end[129][3]) || (phase_count[4] ^ phase_end[129][4]) || (phase_count[5] ^ phase_end[129][5]) || (phase_count[6] ^ phase_end[129][6]) || phase[129][7];
	assign select_end[130] = (phase_count[0] ^ phase_end[130][0]) || (phase_count[1] ^ phase_end[130][1]) || (phase_count[2] ^ phase_end[130][2]) || (phase_count[3] ^ phase_end[130][3]) || (phase_count[4] ^ phase_end[130][4]) || (phase_count[5] ^ phase_end[130][5]) || (phase_count[6] ^ phase_end[130][6]) || phase[130][7];
	assign select_end[131] = (phase_count[0] ^ phase_end[131][0]) || (phase_count[1] ^ phase_end[131][1]) || (phase_count[2] ^ phase_end[131][2]) || (phase_count[3] ^ phase_end[131][3]) || (phase_count[4] ^ phase_end[131][4]) || (phase_count[5] ^ phase_end[131][5]) || (phase_count[6] ^ phase_end[131][6]) || phase[131][7];
	assign select_end[132] = (phase_count[0] ^ phase_end[132][0]) || (phase_count[1] ^ phase_end[132][1]) || (phase_count[2] ^ phase_end[132][2]) || (phase_count[3] ^ phase_end[132][3]) || (phase_count[4] ^ phase_end[132][4]) || (phase_count[5] ^ phase_end[132][5]) || (phase_count[6] ^ phase_end[132][6]) || phase[132][7];
	assign select_end[133] = (phase_count[0] ^ phase_end[133][0]) || (phase_count[1] ^ phase_end[133][1]) || (phase_count[2] ^ phase_end[133][2]) || (phase_count[3] ^ phase_end[133][3]) || (phase_count[4] ^ phase_end[133][4]) || (phase_count[5] ^ phase_end[133][5]) || (phase_count[6] ^ phase_end[133][6]) || phase[133][7];
	assign select_end[134] = (phase_count[0] ^ phase_end[134][0]) || (phase_count[1] ^ phase_end[134][1]) || (phase_count[2] ^ phase_end[134][2]) || (phase_count[3] ^ phase_end[134][3]) || (phase_count[4] ^ phase_end[134][4]) || (phase_count[5] ^ phase_end[134][5]) || (phase_count[6] ^ phase_end[134][6]) || phase[134][7];
	assign select_end[135] = (phase_count[0] ^ phase_end[135][0]) || (phase_count[1] ^ phase_end[135][1]) || (phase_count[2] ^ phase_end[135][2]) || (phase_count[3] ^ phase_end[135][3]) || (phase_count[4] ^ phase_end[135][4]) || (phase_count[5] ^ phase_end[135][5]) || (phase_count[6] ^ phase_end[135][6]) || phase[135][7];
	assign select_end[136] = (phase_count[0] ^ phase_end[136][0]) || (phase_count[1] ^ phase_end[136][1]) || (phase_count[2] ^ phase_end[136][2]) || (phase_count[3] ^ phase_end[136][3]) || (phase_count[4] ^ phase_end[136][4]) || (phase_count[5] ^ phase_end[136][5]) || (phase_count[6] ^ phase_end[136][6]) || phase[136][7];
	assign select_end[137] = (phase_count[0] ^ phase_end[137][0]) || (phase_count[1] ^ phase_end[137][1]) || (phase_count[2] ^ phase_end[137][2]) || (phase_count[3] ^ phase_end[137][3]) || (phase_count[4] ^ phase_end[137][4]) || (phase_count[5] ^ phase_end[137][5]) || (phase_count[6] ^ phase_end[137][6]) || phase[137][7];
	assign select_end[138] = (phase_count[0] ^ phase_end[138][0]) || (phase_count[1] ^ phase_end[138][1]) || (phase_count[2] ^ phase_end[138][2]) || (phase_count[3] ^ phase_end[138][3]) || (phase_count[4] ^ phase_end[138][4]) || (phase_count[5] ^ phase_end[138][5]) || (phase_count[6] ^ phase_end[138][6]) || phase[138][7];
	assign select_end[139] = (phase_count[0] ^ phase_end[139][0]) || (phase_count[1] ^ phase_end[139][1]) || (phase_count[2] ^ phase_end[139][2]) || (phase_count[3] ^ phase_end[139][3]) || (phase_count[4] ^ phase_end[139][4]) || (phase_count[5] ^ phase_end[139][5]) || (phase_count[6] ^ phase_end[139][6]) || phase[139][7];
	assign select_end[140] = (phase_count[0] ^ phase_end[140][0]) || (phase_count[1] ^ phase_end[140][1]) || (phase_count[2] ^ phase_end[140][2]) || (phase_count[3] ^ phase_end[140][3]) || (phase_count[4] ^ phase_end[140][4]) || (phase_count[5] ^ phase_end[140][5]) || (phase_count[6] ^ phase_end[140][6]) || phase[140][7];
	assign select_end[141] = (phase_count[0] ^ phase_end[141][0]) || (phase_count[1] ^ phase_end[141][1]) || (phase_count[2] ^ phase_end[141][2]) || (phase_count[3] ^ phase_end[141][3]) || (phase_count[4] ^ phase_end[141][4]) || (phase_count[5] ^ phase_end[141][5]) || (phase_count[6] ^ phase_end[141][6]) || phase[141][7];
	assign select_end[142] = (phase_count[0] ^ phase_end[142][0]) || (phase_count[1] ^ phase_end[142][1]) || (phase_count[2] ^ phase_end[142][2]) || (phase_count[3] ^ phase_end[142][3]) || (phase_count[4] ^ phase_end[142][4]) || (phase_count[5] ^ phase_end[142][5]) || (phase_count[6] ^ phase_end[142][6]) || phase[142][7];
	assign select_end[143] = (phase_count[0] ^ phase_end[143][0]) || (phase_count[1] ^ phase_end[143][1]) || (phase_count[2] ^ phase_end[143][2]) || (phase_count[3] ^ phase_end[143][3]) || (phase_count[4] ^ phase_end[143][4]) || (phase_count[5] ^ phase_end[143][5]) || (phase_count[6] ^ phase_end[143][6]) || phase[143][7];
	assign select_end[144] = (phase_count[0] ^ phase_end[144][0]) || (phase_count[1] ^ phase_end[144][1]) || (phase_count[2] ^ phase_end[144][2]) || (phase_count[3] ^ phase_end[144][3]) || (phase_count[4] ^ phase_end[144][4]) || (phase_count[5] ^ phase_end[144][5]) || (phase_count[6] ^ phase_end[144][6]) || phase[144][7];
	assign select_end[145] = (phase_count[0] ^ phase_end[145][0]) || (phase_count[1] ^ phase_end[145][1]) || (phase_count[2] ^ phase_end[145][2]) || (phase_count[3] ^ phase_end[145][3]) || (phase_count[4] ^ phase_end[145][4]) || (phase_count[5] ^ phase_end[145][5]) || (phase_count[6] ^ phase_end[145][6]) || phase[145][7];
	assign select_end[146] = (phase_count[0] ^ phase_end[146][0]) || (phase_count[1] ^ phase_end[146][1]) || (phase_count[2] ^ phase_end[146][2]) || (phase_count[3] ^ phase_end[146][3]) || (phase_count[4] ^ phase_end[146][4]) || (phase_count[5] ^ phase_end[146][5]) || (phase_count[6] ^ phase_end[146][6]) || phase[146][7];
	assign select_end[147] = (phase_count[0] ^ phase_end[147][0]) || (phase_count[1] ^ phase_end[147][1]) || (phase_count[2] ^ phase_end[147][2]) || (phase_count[3] ^ phase_end[147][3]) || (phase_count[4] ^ phase_end[147][4]) || (phase_count[5] ^ phase_end[147][5]) || (phase_count[6] ^ phase_end[147][6]) || phase[147][7];
	assign select_end[148] = (phase_count[0] ^ phase_end[148][0]) || (phase_count[1] ^ phase_end[148][1]) || (phase_count[2] ^ phase_end[148][2]) || (phase_count[3] ^ phase_end[148][3]) || (phase_count[4] ^ phase_end[148][4]) || (phase_count[5] ^ phase_end[148][5]) || (phase_count[6] ^ phase_end[148][6]) || phase[148][7];
	assign select_end[149] = (phase_count[0] ^ phase_end[149][0]) || (phase_count[1] ^ phase_end[149][1]) || (phase_count[2] ^ phase_end[149][2]) || (phase_count[3] ^ phase_end[149][3]) || (phase_count[4] ^ phase_end[149][4]) || (phase_count[5] ^ phase_end[149][5]) || (phase_count[6] ^ phase_end[149][6]) || phase[149][7];
	assign select_end[150] = (phase_count[0] ^ phase_end[150][0]) || (phase_count[1] ^ phase_end[150][1]) || (phase_count[2] ^ phase_end[150][2]) || (phase_count[3] ^ phase_end[150][3]) || (phase_count[4] ^ phase_end[150][4]) || (phase_count[5] ^ phase_end[150][5]) || (phase_count[6] ^ phase_end[150][6]) || phase[150][7];
	assign select_end[151] = (phase_count[0] ^ phase_end[151][0]) || (phase_count[1] ^ phase_end[151][1]) || (phase_count[2] ^ phase_end[151][2]) || (phase_count[3] ^ phase_end[151][3]) || (phase_count[4] ^ phase_end[151][4]) || (phase_count[5] ^ phase_end[151][5]) || (phase_count[6] ^ phase_end[151][6]) || phase[151][7];
	assign select_end[152] = (phase_count[0] ^ phase_end[152][0]) || (phase_count[1] ^ phase_end[152][1]) || (phase_count[2] ^ phase_end[152][2]) || (phase_count[3] ^ phase_end[152][3]) || (phase_count[4] ^ phase_end[152][4]) || (phase_count[5] ^ phase_end[152][5]) || (phase_count[6] ^ phase_end[152][6]) || phase[152][7];
	assign select_end[153] = (phase_count[0] ^ phase_end[153][0]) || (phase_count[1] ^ phase_end[153][1]) || (phase_count[2] ^ phase_end[153][2]) || (phase_count[3] ^ phase_end[153][3]) || (phase_count[4] ^ phase_end[153][4]) || (phase_count[5] ^ phase_end[153][5]) || (phase_count[6] ^ phase_end[153][6]) || phase[153][7];
	assign select_end[154] = (phase_count[0] ^ phase_end[154][0]) || (phase_count[1] ^ phase_end[154][1]) || (phase_count[2] ^ phase_end[154][2]) || (phase_count[3] ^ phase_end[154][3]) || (phase_count[4] ^ phase_end[154][4]) || (phase_count[5] ^ phase_end[154][5]) || (phase_count[6] ^ phase_end[154][6]) || phase[154][7];
	assign select_end[155] = (phase_count[0] ^ phase_end[155][0]) || (phase_count[1] ^ phase_end[155][1]) || (phase_count[2] ^ phase_end[155][2]) || (phase_count[3] ^ phase_end[155][3]) || (phase_count[4] ^ phase_end[155][4]) || (phase_count[5] ^ phase_end[155][5]) || (phase_count[6] ^ phase_end[155][6]) || phase[155][7];
	assign select_end[156] = (phase_count[0] ^ phase_end[156][0]) || (phase_count[1] ^ phase_end[156][1]) || (phase_count[2] ^ phase_end[156][2]) || (phase_count[3] ^ phase_end[156][3]) || (phase_count[4] ^ phase_end[156][4]) || (phase_count[5] ^ phase_end[156][5]) || (phase_count[6] ^ phase_end[156][6]) || phase[156][7];
	assign select_end[157] = (phase_count[0] ^ phase_end[157][0]) || (phase_count[1] ^ phase_end[157][1]) || (phase_count[2] ^ phase_end[157][2]) || (phase_count[3] ^ phase_end[157][3]) || (phase_count[4] ^ phase_end[157][4]) || (phase_count[5] ^ phase_end[157][5]) || (phase_count[6] ^ phase_end[157][6]) || phase[157][7];
	assign select_end[158] = (phase_count[0] ^ phase_end[158][0]) || (phase_count[1] ^ phase_end[158][1]) || (phase_count[2] ^ phase_end[158][2]) || (phase_count[3] ^ phase_end[158][3]) || (phase_count[4] ^ phase_end[158][4]) || (phase_count[5] ^ phase_end[158][5]) || (phase_count[6] ^ phase_end[158][6]) || phase[158][7];
	assign select_end[159] = (phase_count[0] ^ phase_end[159][0]) || (phase_count[1] ^ phase_end[159][1]) || (phase_count[2] ^ phase_end[159][2]) || (phase_count[3] ^ phase_end[159][3]) || (phase_count[4] ^ phase_end[159][4]) || (phase_count[5] ^ phase_end[159][5]) || (phase_count[6] ^ phase_end[159][6]) || phase[159][7];
	assign select_end[160] = (phase_count[0] ^ phase_end[160][0]) || (phase_count[1] ^ phase_end[160][1]) || (phase_count[2] ^ phase_end[160][2]) || (phase_count[3] ^ phase_end[160][3]) || (phase_count[4] ^ phase_end[160][4]) || (phase_count[5] ^ phase_end[160][5]) || (phase_count[6] ^ phase_end[160][6]) || phase[160][7];
	assign select_end[161] = (phase_count[0] ^ phase_end[161][0]) || (phase_count[1] ^ phase_end[161][1]) || (phase_count[2] ^ phase_end[161][2]) || (phase_count[3] ^ phase_end[161][3]) || (phase_count[4] ^ phase_end[161][4]) || (phase_count[5] ^ phase_end[161][5]) || (phase_count[6] ^ phase_end[161][6]) || phase[161][7];
	assign select_end[162] = (phase_count[0] ^ phase_end[162][0]) || (phase_count[1] ^ phase_end[162][1]) || (phase_count[2] ^ phase_end[162][2]) || (phase_count[3] ^ phase_end[162][3]) || (phase_count[4] ^ phase_end[162][4]) || (phase_count[5] ^ phase_end[162][5]) || (phase_count[6] ^ phase_end[162][6]) || phase[162][7];
	assign select_end[163] = (phase_count[0] ^ phase_end[163][0]) || (phase_count[1] ^ phase_end[163][1]) || (phase_count[2] ^ phase_end[163][2]) || (phase_count[3] ^ phase_end[163][3]) || (phase_count[4] ^ phase_end[163][4]) || (phase_count[5] ^ phase_end[163][5]) || (phase_count[6] ^ phase_end[163][6]) || phase[163][7];
	assign select_end[164] = (phase_count[0] ^ phase_end[164][0]) || (phase_count[1] ^ phase_end[164][1]) || (phase_count[2] ^ phase_end[164][2]) || (phase_count[3] ^ phase_end[164][3]) || (phase_count[4] ^ phase_end[164][4]) || (phase_count[5] ^ phase_end[164][5]) || (phase_count[6] ^ phase_end[164][6]) || phase[164][7];
	assign select_end[165] = (phase_count[0] ^ phase_end[165][0]) || (phase_count[1] ^ phase_end[165][1]) || (phase_count[2] ^ phase_end[165][2]) || (phase_count[3] ^ phase_end[165][3]) || (phase_count[4] ^ phase_end[165][4]) || (phase_count[5] ^ phase_end[165][5]) || (phase_count[6] ^ phase_end[165][6]) || phase[165][7];
	assign select_end[166] = (phase_count[0] ^ phase_end[166][0]) || (phase_count[1] ^ phase_end[166][1]) || (phase_count[2] ^ phase_end[166][2]) || (phase_count[3] ^ phase_end[166][3]) || (phase_count[4] ^ phase_end[166][4]) || (phase_count[5] ^ phase_end[166][5]) || (phase_count[6] ^ phase_end[166][6]) || phase[166][7];
	assign select_end[167] = (phase_count[0] ^ phase_end[167][0]) || (phase_count[1] ^ phase_end[167][1]) || (phase_count[2] ^ phase_end[167][2]) || (phase_count[3] ^ phase_end[167][3]) || (phase_count[4] ^ phase_end[167][4]) || (phase_count[5] ^ phase_end[167][5]) || (phase_count[6] ^ phase_end[167][6]) || phase[167][7];
	assign select_end[168] = (phase_count[0] ^ phase_end[168][0]) || (phase_count[1] ^ phase_end[168][1]) || (phase_count[2] ^ phase_end[168][2]) || (phase_count[3] ^ phase_end[168][3]) || (phase_count[4] ^ phase_end[168][4]) || (phase_count[5] ^ phase_end[168][5]) || (phase_count[6] ^ phase_end[168][6]) || phase[168][7];
	assign select_end[169] = (phase_count[0] ^ phase_end[169][0]) || (phase_count[1] ^ phase_end[169][1]) || (phase_count[2] ^ phase_end[169][2]) || (phase_count[3] ^ phase_end[169][3]) || (phase_count[4] ^ phase_end[169][4]) || (phase_count[5] ^ phase_end[169][5]) || (phase_count[6] ^ phase_end[169][6]) || phase[169][7];
	assign select_end[170] = (phase_count[0] ^ phase_end[170][0]) || (phase_count[1] ^ phase_end[170][1]) || (phase_count[2] ^ phase_end[170][2]) || (phase_count[3] ^ phase_end[170][3]) || (phase_count[4] ^ phase_end[170][4]) || (phase_count[5] ^ phase_end[170][5]) || (phase_count[6] ^ phase_end[170][6]) || phase[170][7];
	assign select_end[171] = (phase_count[0] ^ phase_end[171][0]) || (phase_count[1] ^ phase_end[171][1]) || (phase_count[2] ^ phase_end[171][2]) || (phase_count[3] ^ phase_end[171][3]) || (phase_count[4] ^ phase_end[171][4]) || (phase_count[5] ^ phase_end[171][5]) || (phase_count[6] ^ phase_end[171][6]) || phase[171][7];
	assign select_end[172] = (phase_count[0] ^ phase_end[172][0]) || (phase_count[1] ^ phase_end[172][1]) || (phase_count[2] ^ phase_end[172][2]) || (phase_count[3] ^ phase_end[172][3]) || (phase_count[4] ^ phase_end[172][4]) || (phase_count[5] ^ phase_end[172][5]) || (phase_count[6] ^ phase_end[172][6]) || phase[172][7];
	assign select_end[173] = (phase_count[0] ^ phase_end[173][0]) || (phase_count[1] ^ phase_end[173][1]) || (phase_count[2] ^ phase_end[173][2]) || (phase_count[3] ^ phase_end[173][3]) || (phase_count[4] ^ phase_end[173][4]) || (phase_count[5] ^ phase_end[173][5]) || (phase_count[6] ^ phase_end[173][6]) || phase[173][7];
	assign select_end[174] = (phase_count[0] ^ phase_end[174][0]) || (phase_count[1] ^ phase_end[174][1]) || (phase_count[2] ^ phase_end[174][2]) || (phase_count[3] ^ phase_end[174][3]) || (phase_count[4] ^ phase_end[174][4]) || (phase_count[5] ^ phase_end[174][5]) || (phase_count[6] ^ phase_end[174][6]) || phase[174][7];
	assign select_end[175] = (phase_count[0] ^ phase_end[175][0]) || (phase_count[1] ^ phase_end[175][1]) || (phase_count[2] ^ phase_end[175][2]) || (phase_count[3] ^ phase_end[175][3]) || (phase_count[4] ^ phase_end[175][4]) || (phase_count[5] ^ phase_end[175][5]) || (phase_count[6] ^ phase_end[175][6]) || phase[175][7];
	assign select_end[176] = (phase_count[0] ^ phase_end[176][0]) || (phase_count[1] ^ phase_end[176][1]) || (phase_count[2] ^ phase_end[176][2]) || (phase_count[3] ^ phase_end[176][3]) || (phase_count[4] ^ phase_end[176][4]) || (phase_count[5] ^ phase_end[176][5]) || (phase_count[6] ^ phase_end[176][6]) || phase[176][7];
	assign select_end[177] = (phase_count[0] ^ phase_end[177][0]) || (phase_count[1] ^ phase_end[177][1]) || (phase_count[2] ^ phase_end[177][2]) || (phase_count[3] ^ phase_end[177][3]) || (phase_count[4] ^ phase_end[177][4]) || (phase_count[5] ^ phase_end[177][5]) || (phase_count[6] ^ phase_end[177][6]) || phase[177][7];
	assign select_end[178] = (phase_count[0] ^ phase_end[178][0]) || (phase_count[1] ^ phase_end[178][1]) || (phase_count[2] ^ phase_end[178][2]) || (phase_count[3] ^ phase_end[178][3]) || (phase_count[4] ^ phase_end[178][4]) || (phase_count[5] ^ phase_end[178][5]) || (phase_count[6] ^ phase_end[178][6]) || phase[178][7];
	assign select_end[179] = (phase_count[0] ^ phase_end[179][0]) || (phase_count[1] ^ phase_end[179][1]) || (phase_count[2] ^ phase_end[179][2]) || (phase_count[3] ^ phase_end[179][3]) || (phase_count[4] ^ phase_end[179][4]) || (phase_count[5] ^ phase_end[179][5]) || (phase_count[6] ^ phase_end[179][6]) || phase[179][7];
	assign select_end[180] = (phase_count[0] ^ phase_end[180][0]) || (phase_count[1] ^ phase_end[180][1]) || (phase_count[2] ^ phase_end[180][2]) || (phase_count[3] ^ phase_end[180][3]) || (phase_count[4] ^ phase_end[180][4]) || (phase_count[5] ^ phase_end[180][5]) || (phase_count[6] ^ phase_end[180][6]) || phase[180][7];
	assign select_end[181] = (phase_count[0] ^ phase_end[181][0]) || (phase_count[1] ^ phase_end[181][1]) || (phase_count[2] ^ phase_end[181][2]) || (phase_count[3] ^ phase_end[181][3]) || (phase_count[4] ^ phase_end[181][4]) || (phase_count[5] ^ phase_end[181][5]) || (phase_count[6] ^ phase_end[181][6]) || phase[181][7];
	assign select_end[182] = (phase_count[0] ^ phase_end[182][0]) || (phase_count[1] ^ phase_end[182][1]) || (phase_count[2] ^ phase_end[182][2]) || (phase_count[3] ^ phase_end[182][3]) || (phase_count[4] ^ phase_end[182][4]) || (phase_count[5] ^ phase_end[182][5]) || (phase_count[6] ^ phase_end[182][6]) || phase[182][7];
	assign select_end[183] = (phase_count[0] ^ phase_end[183][0]) || (phase_count[1] ^ phase_end[183][1]) || (phase_count[2] ^ phase_end[183][2]) || (phase_count[3] ^ phase_end[183][3]) || (phase_count[4] ^ phase_end[183][4]) || (phase_count[5] ^ phase_end[183][5]) || (phase_count[6] ^ phase_end[183][6]) || phase[183][7];
	assign select_end[184] = (phase_count[0] ^ phase_end[184][0]) || (phase_count[1] ^ phase_end[184][1]) || (phase_count[2] ^ phase_end[184][2]) || (phase_count[3] ^ phase_end[184][3]) || (phase_count[4] ^ phase_end[184][4]) || (phase_count[5] ^ phase_end[184][5]) || (phase_count[6] ^ phase_end[184][6]) || phase[184][7];
	assign select_end[185] = (phase_count[0] ^ phase_end[185][0]) || (phase_count[1] ^ phase_end[185][1]) || (phase_count[2] ^ phase_end[185][2]) || (phase_count[3] ^ phase_end[185][3]) || (phase_count[4] ^ phase_end[185][4]) || (phase_count[5] ^ phase_end[185][5]) || (phase_count[6] ^ phase_end[185][6]) || phase[185][7];
	assign select_end[186] = (phase_count[0] ^ phase_end[186][0]) || (phase_count[1] ^ phase_end[186][1]) || (phase_count[2] ^ phase_end[186][2]) || (phase_count[3] ^ phase_end[186][3]) || (phase_count[4] ^ phase_end[186][4]) || (phase_count[5] ^ phase_end[186][5]) || (phase_count[6] ^ phase_end[186][6]) || phase[186][7];
	assign select_end[187] = (phase_count[0] ^ phase_end[187][0]) || (phase_count[1] ^ phase_end[187][1]) || (phase_count[2] ^ phase_end[187][2]) || (phase_count[3] ^ phase_end[187][3]) || (phase_count[4] ^ phase_end[187][4]) || (phase_count[5] ^ phase_end[187][5]) || (phase_count[6] ^ phase_end[187][6]) || phase[187][7];
	assign select_end[188] = (phase_count[0] ^ phase_end[188][0]) || (phase_count[1] ^ phase_end[188][1]) || (phase_count[2] ^ phase_end[188][2]) || (phase_count[3] ^ phase_end[188][3]) || (phase_count[4] ^ phase_end[188][4]) || (phase_count[5] ^ phase_end[188][5]) || (phase_count[6] ^ phase_end[188][6]) || phase[188][7];
	assign select_end[189] = (phase_count[0] ^ phase_end[189][0]) || (phase_count[1] ^ phase_end[189][1]) || (phase_count[2] ^ phase_end[189][2]) || (phase_count[3] ^ phase_end[189][3]) || (phase_count[4] ^ phase_end[189][4]) || (phase_count[5] ^ phase_end[189][5]) || (phase_count[6] ^ phase_end[189][6]) || phase[189][7];
	assign select_end[190] = (phase_count[0] ^ phase_end[190][0]) || (phase_count[1] ^ phase_end[190][1]) || (phase_count[2] ^ phase_end[190][2]) || (phase_count[3] ^ phase_end[190][3]) || (phase_count[4] ^ phase_end[190][4]) || (phase_count[5] ^ phase_end[190][5]) || (phase_count[6] ^ phase_end[190][6]) || phase[190][7];
	assign select_end[191] = (phase_count[0] ^ phase_end[191][0]) || (phase_count[1] ^ phase_end[191][1]) || (phase_count[2] ^ phase_end[191][2]) || (phase_count[3] ^ phase_end[191][3]) || (phase_count[4] ^ phase_end[191][4]) || (phase_count[5] ^ phase_end[191][5]) || (phase_count[6] ^ phase_end[191][6]) || phase[191][7];
	assign select_end[192] = (phase_count[0] ^ phase_end[192][0]) || (phase_count[1] ^ phase_end[192][1]) || (phase_count[2] ^ phase_end[192][2]) || (phase_count[3] ^ phase_end[192][3]) || (phase_count[4] ^ phase_end[192][4]) || (phase_count[5] ^ phase_end[192][5]) || (phase_count[6] ^ phase_end[192][6]) || phase[192][7];
	assign select_end[193] = (phase_count[0] ^ phase_end[193][0]) || (phase_count[1] ^ phase_end[193][1]) || (phase_count[2] ^ phase_end[193][2]) || (phase_count[3] ^ phase_end[193][3]) || (phase_count[4] ^ phase_end[193][4]) || (phase_count[5] ^ phase_end[193][5]) || (phase_count[6] ^ phase_end[193][6]) || phase[193][7];
	assign select_end[194] = (phase_count[0] ^ phase_end[194][0]) || (phase_count[1] ^ phase_end[194][1]) || (phase_count[2] ^ phase_end[194][2]) || (phase_count[3] ^ phase_end[194][3]) || (phase_count[4] ^ phase_end[194][4]) || (phase_count[5] ^ phase_end[194][5]) || (phase_count[6] ^ phase_end[194][6]) || phase[194][7];
	assign select_end[195] = (phase_count[0] ^ phase_end[195][0]) || (phase_count[1] ^ phase_end[195][1]) || (phase_count[2] ^ phase_end[195][2]) || (phase_count[3] ^ phase_end[195][3]) || (phase_count[4] ^ phase_end[195][4]) || (phase_count[5] ^ phase_end[195][5]) || (phase_count[6] ^ phase_end[195][6]) || phase[195][7];
	assign select_end[196] = (phase_count[0] ^ phase_end[196][0]) || (phase_count[1] ^ phase_end[196][1]) || (phase_count[2] ^ phase_end[196][2]) || (phase_count[3] ^ phase_end[196][3]) || (phase_count[4] ^ phase_end[196][4]) || (phase_count[5] ^ phase_end[196][5]) || (phase_count[6] ^ phase_end[196][6]) || phase[196][7];
	assign select_end[197] = (phase_count[0] ^ phase_end[197][0]) || (phase_count[1] ^ phase_end[197][1]) || (phase_count[2] ^ phase_end[197][2]) || (phase_count[3] ^ phase_end[197][3]) || (phase_count[4] ^ phase_end[197][4]) || (phase_count[5] ^ phase_end[197][5]) || (phase_count[6] ^ phase_end[197][6]) || phase[197][7];
	assign select_end[198] = (phase_count[0] ^ phase_end[198][0]) || (phase_count[1] ^ phase_end[198][1]) || (phase_count[2] ^ phase_end[198][2]) || (phase_count[3] ^ phase_end[198][3]) || (phase_count[4] ^ phase_end[198][4]) || (phase_count[5] ^ phase_end[198][5]) || (phase_count[6] ^ phase_end[198][6]) || phase[198][7];
	assign select_end[199] = (phase_count[0] ^ phase_end[199][0]) || (phase_count[1] ^ phase_end[199][1]) || (phase_count[2] ^ phase_end[199][2]) || (phase_count[3] ^ phase_end[199][3]) || (phase_count[4] ^ phase_end[199][4]) || (phase_count[5] ^ phase_end[199][5]) || (phase_count[6] ^ phase_end[199][6]) || phase[199][7];
	assign select_end[200] = (phase_count[0] ^ phase_end[200][0]) || (phase_count[1] ^ phase_end[200][1]) || (phase_count[2] ^ phase_end[200][2]) || (phase_count[3] ^ phase_end[200][3]) || (phase_count[4] ^ phase_end[200][4]) || (phase_count[5] ^ phase_end[200][5]) || (phase_count[6] ^ phase_end[200][6]) || phase[200][7];
	assign select_end[201] = (phase_count[0] ^ phase_end[201][0]) || (phase_count[1] ^ phase_end[201][1]) || (phase_count[2] ^ phase_end[201][2]) || (phase_count[3] ^ phase_end[201][3]) || (phase_count[4] ^ phase_end[201][4]) || (phase_count[5] ^ phase_end[201][5]) || (phase_count[6] ^ phase_end[201][6]) || phase[201][7];
	assign select_end[202] = (phase_count[0] ^ phase_end[202][0]) || (phase_count[1] ^ phase_end[202][1]) || (phase_count[2] ^ phase_end[202][2]) || (phase_count[3] ^ phase_end[202][3]) || (phase_count[4] ^ phase_end[202][4]) || (phase_count[5] ^ phase_end[202][5]) || (phase_count[6] ^ phase_end[202][6]) || phase[202][7];
	assign select_end[203] = (phase_count[0] ^ phase_end[203][0]) || (phase_count[1] ^ phase_end[203][1]) || (phase_count[2] ^ phase_end[203][2]) || (phase_count[3] ^ phase_end[203][3]) || (phase_count[4] ^ phase_end[203][4]) || (phase_count[5] ^ phase_end[203][5]) || (phase_count[6] ^ phase_end[203][6]) || phase[203][7];
	assign select_end[204] = (phase_count[0] ^ phase_end[204][0]) || (phase_count[1] ^ phase_end[204][1]) || (phase_count[2] ^ phase_end[204][2]) || (phase_count[3] ^ phase_end[204][3]) || (phase_count[4] ^ phase_end[204][4]) || (phase_count[5] ^ phase_end[204][5]) || (phase_count[6] ^ phase_end[204][6]) || phase[204][7];
	assign select_end[205] = (phase_count[0] ^ phase_end[205][0]) || (phase_count[1] ^ phase_end[205][1]) || (phase_count[2] ^ phase_end[205][2]) || (phase_count[3] ^ phase_end[205][3]) || (phase_count[4] ^ phase_end[205][4]) || (phase_count[5] ^ phase_end[205][5]) || (phase_count[6] ^ phase_end[205][6]) || phase[205][7];
	assign select_end[206] = (phase_count[0] ^ phase_end[206][0]) || (phase_count[1] ^ phase_end[206][1]) || (phase_count[2] ^ phase_end[206][2]) || (phase_count[3] ^ phase_end[206][3]) || (phase_count[4] ^ phase_end[206][4]) || (phase_count[5] ^ phase_end[206][5]) || (phase_count[6] ^ phase_end[206][6]) || phase[206][7];
	assign select_end[207] = (phase_count[0] ^ phase_end[207][0]) || (phase_count[1] ^ phase_end[207][1]) || (phase_count[2] ^ phase_end[207][2]) || (phase_count[3] ^ phase_end[207][3]) || (phase_count[4] ^ phase_end[207][4]) || (phase_count[5] ^ phase_end[207][5]) || (phase_count[6] ^ phase_end[207][6]) || phase[207][7];
	assign select_end[208] = (phase_count[0] ^ phase_end[208][0]) || (phase_count[1] ^ phase_end[208][1]) || (phase_count[2] ^ phase_end[208][2]) || (phase_count[3] ^ phase_end[208][3]) || (phase_count[4] ^ phase_end[208][4]) || (phase_count[5] ^ phase_end[208][5]) || (phase_count[6] ^ phase_end[208][6]) || phase[208][7];
	assign select_end[209] = (phase_count[0] ^ phase_end[209][0]) || (phase_count[1] ^ phase_end[209][1]) || (phase_count[2] ^ phase_end[209][2]) || (phase_count[3] ^ phase_end[209][3]) || (phase_count[4] ^ phase_end[209][4]) || (phase_count[5] ^ phase_end[209][5]) || (phase_count[6] ^ phase_end[209][6]) || phase[209][7];
	assign select_end[210] = (phase_count[0] ^ phase_end[210][0]) || (phase_count[1] ^ phase_end[210][1]) || (phase_count[2] ^ phase_end[210][2]) || (phase_count[3] ^ phase_end[210][3]) || (phase_count[4] ^ phase_end[210][4]) || (phase_count[5] ^ phase_end[210][5]) || (phase_count[6] ^ phase_end[210][6]) || phase[210][7];
	assign select_end[211] = (phase_count[0] ^ phase_end[211][0]) || (phase_count[1] ^ phase_end[211][1]) || (phase_count[2] ^ phase_end[211][2]) || (phase_count[3] ^ phase_end[211][3]) || (phase_count[4] ^ phase_end[211][4]) || (phase_count[5] ^ phase_end[211][5]) || (phase_count[6] ^ phase_end[211][6]) || phase[211][7];
	assign select_end[212] = (phase_count[0] ^ phase_end[212][0]) || (phase_count[1] ^ phase_end[212][1]) || (phase_count[2] ^ phase_end[212][2]) || (phase_count[3] ^ phase_end[212][3]) || (phase_count[4] ^ phase_end[212][4]) || (phase_count[5] ^ phase_end[212][5]) || (phase_count[6] ^ phase_end[212][6]) || phase[212][7];
	assign select_end[213] = (phase_count[0] ^ phase_end[213][0]) || (phase_count[1] ^ phase_end[213][1]) || (phase_count[2] ^ phase_end[213][2]) || (phase_count[3] ^ phase_end[213][3]) || (phase_count[4] ^ phase_end[213][4]) || (phase_count[5] ^ phase_end[213][5]) || (phase_count[6] ^ phase_end[213][6]) || phase[213][7];
	assign select_end[214] = (phase_count[0] ^ phase_end[214][0]) || (phase_count[1] ^ phase_end[214][1]) || (phase_count[2] ^ phase_end[214][2]) || (phase_count[3] ^ phase_end[214][3]) || (phase_count[4] ^ phase_end[214][4]) || (phase_count[5] ^ phase_end[214][5]) || (phase_count[6] ^ phase_end[214][6]) || phase[214][7];
	assign select_end[215] = (phase_count[0] ^ phase_end[215][0]) || (phase_count[1] ^ phase_end[215][1]) || (phase_count[2] ^ phase_end[215][2]) || (phase_count[3] ^ phase_end[215][3]) || (phase_count[4] ^ phase_end[215][4]) || (phase_count[5] ^ phase_end[215][5]) || (phase_count[6] ^ phase_end[215][6]) || phase[215][7];
	assign select_end[216] = (phase_count[0] ^ phase_end[216][0]) || (phase_count[1] ^ phase_end[216][1]) || (phase_count[2] ^ phase_end[216][2]) || (phase_count[3] ^ phase_end[216][3]) || (phase_count[4] ^ phase_end[216][4]) || (phase_count[5] ^ phase_end[216][5]) || (phase_count[6] ^ phase_end[216][6]) || phase[216][7];
	assign select_end[217] = (phase_count[0] ^ phase_end[217][0]) || (phase_count[1] ^ phase_end[217][1]) || (phase_count[2] ^ phase_end[217][2]) || (phase_count[3] ^ phase_end[217][3]) || (phase_count[4] ^ phase_end[217][4]) || (phase_count[5] ^ phase_end[217][5]) || (phase_count[6] ^ phase_end[217][6]) || phase[217][7];
	assign select_end[218] = (phase_count[0] ^ phase_end[218][0]) || (phase_count[1] ^ phase_end[218][1]) || (phase_count[2] ^ phase_end[218][2]) || (phase_count[3] ^ phase_end[218][3]) || (phase_count[4] ^ phase_end[218][4]) || (phase_count[5] ^ phase_end[218][5]) || (phase_count[6] ^ phase_end[218][6]) || phase[218][7];
	assign select_end[219] = (phase_count[0] ^ phase_end[219][0]) || (phase_count[1] ^ phase_end[219][1]) || (phase_count[2] ^ phase_end[219][2]) || (phase_count[3] ^ phase_end[219][3]) || (phase_count[4] ^ phase_end[219][4]) || (phase_count[5] ^ phase_end[219][5]) || (phase_count[6] ^ phase_end[219][6]) || phase[219][7];
	assign select_end[220] = (phase_count[0] ^ phase_end[220][0]) || (phase_count[1] ^ phase_end[220][1]) || (phase_count[2] ^ phase_end[220][2]) || (phase_count[3] ^ phase_end[220][3]) || (phase_count[4] ^ phase_end[220][4]) || (phase_count[5] ^ phase_end[220][5]) || (phase_count[6] ^ phase_end[220][6]) || phase[220][7];
	assign select_end[221] = (phase_count[0] ^ phase_end[221][0]) || (phase_count[1] ^ phase_end[221][1]) || (phase_count[2] ^ phase_end[221][2]) || (phase_count[3] ^ phase_end[221][3]) || (phase_count[4] ^ phase_end[221][4]) || (phase_count[5] ^ phase_end[221][5]) || (phase_count[6] ^ phase_end[221][6]) || phase[221][7];
	assign select_end[222] = (phase_count[0] ^ phase_end[222][0]) || (phase_count[1] ^ phase_end[222][1]) || (phase_count[2] ^ phase_end[222][2]) || (phase_count[3] ^ phase_end[222][3]) || (phase_count[4] ^ phase_end[222][4]) || (phase_count[5] ^ phase_end[222][5]) || (phase_count[6] ^ phase_end[222][6]) || phase[222][7];
	assign select_end[223] = (phase_count[0] ^ phase_end[223][0]) || (phase_count[1] ^ phase_end[223][1]) || (phase_count[2] ^ phase_end[223][2]) || (phase_count[3] ^ phase_end[223][3]) || (phase_count[4] ^ phase_end[223][4]) || (phase_count[5] ^ phase_end[223][5]) || (phase_count[6] ^ phase_end[223][6]) || phase[223][7];
	assign select_end[224] = (phase_count[0] ^ phase_end[224][0]) || (phase_count[1] ^ phase_end[224][1]) || (phase_count[2] ^ phase_end[224][2]) || (phase_count[3] ^ phase_end[224][3]) || (phase_count[4] ^ phase_end[224][4]) || (phase_count[5] ^ phase_end[224][5]) || (phase_count[6] ^ phase_end[224][6]) || phase[224][7];
	assign select_end[225] = (phase_count[0] ^ phase_end[225][0]) || (phase_count[1] ^ phase_end[225][1]) || (phase_count[2] ^ phase_end[225][2]) || (phase_count[3] ^ phase_end[225][3]) || (phase_count[4] ^ phase_end[225][4]) || (phase_count[5] ^ phase_end[225][5]) || (phase_count[6] ^ phase_end[225][6]) || phase[225][7];
	assign select_end[226] = (phase_count[0] ^ phase_end[226][0]) || (phase_count[1] ^ phase_end[226][1]) || (phase_count[2] ^ phase_end[226][2]) || (phase_count[3] ^ phase_end[226][3]) || (phase_count[4] ^ phase_end[226][4]) || (phase_count[5] ^ phase_end[226][5]) || (phase_count[6] ^ phase_end[226][6]) || phase[226][7];
	assign select_end[227] = (phase_count[0] ^ phase_end[227][0]) || (phase_count[1] ^ phase_end[227][1]) || (phase_count[2] ^ phase_end[227][2]) || (phase_count[3] ^ phase_end[227][3]) || (phase_count[4] ^ phase_end[227][4]) || (phase_count[5] ^ phase_end[227][5]) || (phase_count[6] ^ phase_end[227][6]) || phase[227][7];
	assign select_end[228] = (phase_count[0] ^ phase_end[228][0]) || (phase_count[1] ^ phase_end[228][1]) || (phase_count[2] ^ phase_end[228][2]) || (phase_count[3] ^ phase_end[228][3]) || (phase_count[4] ^ phase_end[228][4]) || (phase_count[5] ^ phase_end[228][5]) || (phase_count[6] ^ phase_end[228][6]) || phase[228][7];
	assign select_end[229] = (phase_count[0] ^ phase_end[229][0]) || (phase_count[1] ^ phase_end[229][1]) || (phase_count[2] ^ phase_end[229][2]) || (phase_count[3] ^ phase_end[229][3]) || (phase_count[4] ^ phase_end[229][4]) || (phase_count[5] ^ phase_end[229][5]) || (phase_count[6] ^ phase_end[229][6]) || phase[229][7];
	assign select_end[230] = (phase_count[0] ^ phase_end[230][0]) || (phase_count[1] ^ phase_end[230][1]) || (phase_count[2] ^ phase_end[230][2]) || (phase_count[3] ^ phase_end[230][3]) || (phase_count[4] ^ phase_end[230][4]) || (phase_count[5] ^ phase_end[230][5]) || (phase_count[6] ^ phase_end[230][6]) || phase[230][7];
	assign select_end[231] = (phase_count[0] ^ phase_end[231][0]) || (phase_count[1] ^ phase_end[231][1]) || (phase_count[2] ^ phase_end[231][2]) || (phase_count[3] ^ phase_end[231][3]) || (phase_count[4] ^ phase_end[231][4]) || (phase_count[5] ^ phase_end[231][5]) || (phase_count[6] ^ phase_end[231][6]) || phase[231][7];
	assign select_end[232] = (phase_count[0] ^ phase_end[232][0]) || (phase_count[1] ^ phase_end[232][1]) || (phase_count[2] ^ phase_end[232][2]) || (phase_count[3] ^ phase_end[232][3]) || (phase_count[4] ^ phase_end[232][4]) || (phase_count[5] ^ phase_end[232][5]) || (phase_count[6] ^ phase_end[232][6]) || phase[232][7];
	assign select_end[233] = (phase_count[0] ^ phase_end[233][0]) || (phase_count[1] ^ phase_end[233][1]) || (phase_count[2] ^ phase_end[233][2]) || (phase_count[3] ^ phase_end[233][3]) || (phase_count[4] ^ phase_end[233][4]) || (phase_count[5] ^ phase_end[233][5]) || (phase_count[6] ^ phase_end[233][6]) || phase[233][7];
	assign select_end[234] = (phase_count[0] ^ phase_end[234][0]) || (phase_count[1] ^ phase_end[234][1]) || (phase_count[2] ^ phase_end[234][2]) || (phase_count[3] ^ phase_end[234][3]) || (phase_count[4] ^ phase_end[234][4]) || (phase_count[5] ^ phase_end[234][5]) || (phase_count[6] ^ phase_end[234][6]) || phase[234][7];
	assign select_end[235] = (phase_count[0] ^ phase_end[235][0]) || (phase_count[1] ^ phase_end[235][1]) || (phase_count[2] ^ phase_end[235][2]) || (phase_count[3] ^ phase_end[235][3]) || (phase_count[4] ^ phase_end[235][4]) || (phase_count[5] ^ phase_end[235][5]) || (phase_count[6] ^ phase_end[235][6]) || phase[235][7];
	assign select_end[236] = (phase_count[0] ^ phase_end[236][0]) || (phase_count[1] ^ phase_end[236][1]) || (phase_count[2] ^ phase_end[236][2]) || (phase_count[3] ^ phase_end[236][3]) || (phase_count[4] ^ phase_end[236][4]) || (phase_count[5] ^ phase_end[236][5]) || (phase_count[6] ^ phase_end[236][6]) || phase[236][7];
	assign select_end[237] = (phase_count[0] ^ phase_end[237][0]) || (phase_count[1] ^ phase_end[237][1]) || (phase_count[2] ^ phase_end[237][2]) || (phase_count[3] ^ phase_end[237][3]) || (phase_count[4] ^ phase_end[237][4]) || (phase_count[5] ^ phase_end[237][5]) || (phase_count[6] ^ phase_end[237][6]) || phase[237][7];
	assign select_end[238] = (phase_count[0] ^ phase_end[238][0]) || (phase_count[1] ^ phase_end[238][1]) || (phase_count[2] ^ phase_end[238][2]) || (phase_count[3] ^ phase_end[238][3]) || (phase_count[4] ^ phase_end[238][4]) || (phase_count[5] ^ phase_end[238][5]) || (phase_count[6] ^ phase_end[238][6]) || phase[238][7];
	assign select_end[239] = (phase_count[0] ^ phase_end[239][0]) || (phase_count[1] ^ phase_end[239][1]) || (phase_count[2] ^ phase_end[239][2]) || (phase_count[3] ^ phase_end[239][3]) || (phase_count[4] ^ phase_end[239][4]) || (phase_count[5] ^ phase_end[239][5]) || (phase_count[6] ^ phase_end[239][6]) || phase[239][7];
	assign select_end[240] = (phase_count[0] ^ phase_end[240][0]) || (phase_count[1] ^ phase_end[240][1]) || (phase_count[2] ^ phase_end[240][2]) || (phase_count[3] ^ phase_end[240][3]) || (phase_count[4] ^ phase_end[240][4]) || (phase_count[5] ^ phase_end[240][5]) || (phase_count[6] ^ phase_end[240][6]) || phase[240][7];
	assign select_end[241] = (phase_count[0] ^ phase_end[241][0]) || (phase_count[1] ^ phase_end[241][1]) || (phase_count[2] ^ phase_end[241][2]) || (phase_count[3] ^ phase_end[241][3]) || (phase_count[4] ^ phase_end[241][4]) || (phase_count[5] ^ phase_end[241][5]) || (phase_count[6] ^ phase_end[241][6]) || phase[241][7];
	assign select_end[242] = (phase_count[0] ^ phase_end[242][0]) || (phase_count[1] ^ phase_end[242][1]) || (phase_count[2] ^ phase_end[242][2]) || (phase_count[3] ^ phase_end[242][3]) || (phase_count[4] ^ phase_end[242][4]) || (phase_count[5] ^ phase_end[242][5]) || (phase_count[6] ^ phase_end[242][6]) || phase[242][7];
	assign select_end[243] = (phase_count[0] ^ phase_end[243][0]) || (phase_count[1] ^ phase_end[243][1]) || (phase_count[2] ^ phase_end[243][2]) || (phase_count[3] ^ phase_end[243][3]) || (phase_count[4] ^ phase_end[243][4]) || (phase_count[5] ^ phase_end[243][5]) || (phase_count[6] ^ phase_end[243][6]) || phase[243][7];
	assign select_end[244] = (phase_count[0] ^ phase_end[244][0]) || (phase_count[1] ^ phase_end[244][1]) || (phase_count[2] ^ phase_end[244][2]) || (phase_count[3] ^ phase_end[244][3]) || (phase_count[4] ^ phase_end[244][4]) || (phase_count[5] ^ phase_end[244][5]) || (phase_count[6] ^ phase_end[244][6]) || phase[244][7];
	assign select_end[245] = (phase_count[0] ^ phase_end[245][0]) || (phase_count[1] ^ phase_end[245][1]) || (phase_count[2] ^ phase_end[245][2]) || (phase_count[3] ^ phase_end[245][3]) || (phase_count[4] ^ phase_end[245][4]) || (phase_count[5] ^ phase_end[245][5]) || (phase_count[6] ^ phase_end[245][6]) || phase[245][7];
	assign select_end[246] = (phase_count[0] ^ phase_end[246][0]) || (phase_count[1] ^ phase_end[246][1]) || (phase_count[2] ^ phase_end[246][2]) || (phase_count[3] ^ phase_end[246][3]) || (phase_count[4] ^ phase_end[246][4]) || (phase_count[5] ^ phase_end[246][5]) || (phase_count[6] ^ phase_end[246][6]) || phase[246][7];
	assign select_end[247] = (phase_count[0] ^ phase_end[247][0]) || (phase_count[1] ^ phase_end[247][1]) || (phase_count[2] ^ phase_end[247][2]) || (phase_count[3] ^ phase_end[247][3]) || (phase_count[4] ^ phase_end[247][4]) || (phase_count[5] ^ phase_end[247][5]) || (phase_count[6] ^ phase_end[247][6]) || phase[247][7];
	assign select_end[248] = (phase_count[0] ^ phase_end[248][0]) || (phase_count[1] ^ phase_end[248][1]) || (phase_count[2] ^ phase_end[248][2]) || (phase_count[3] ^ phase_end[248][3]) || (phase_count[4] ^ phase_end[248][4]) || (phase_count[5] ^ phase_end[248][5]) || (phase_count[6] ^ phase_end[248][6]) || phase[248][7];
	assign select_end[249] = (phase_count[0] ^ phase_end[249][0]) || (phase_count[1] ^ phase_end[249][1]) || (phase_count[2] ^ phase_end[249][2]) || (phase_count[3] ^ phase_end[249][3]) || (phase_count[4] ^ phase_end[249][4]) || (phase_count[5] ^ phase_end[249][5]) || (phase_count[6] ^ phase_end[249][6]) || phase[249][7];
	assign select_end[250] = (phase_count[0] ^ phase_end[250][0]) || (phase_count[1] ^ phase_end[250][1]) || (phase_count[2] ^ phase_end[250][2]) || (phase_count[3] ^ phase_end[250][3]) || (phase_count[4] ^ phase_end[250][4]) || (phase_count[5] ^ phase_end[250][5]) || (phase_count[6] ^ phase_end[250][6]) || phase[250][7];
	assign select_end[251] = (phase_count[0] ^ phase_end[251][0]) || (phase_count[1] ^ phase_end[251][1]) || (phase_count[2] ^ phase_end[251][2]) || (phase_count[3] ^ phase_end[251][3]) || (phase_count[4] ^ phase_end[251][4]) || (phase_count[5] ^ phase_end[251][5]) || (phase_count[6] ^ phase_end[251][6]) || phase[251][7];
	assign select_end[252] = (phase_count[0] ^ phase_end[252][0]) || (phase_count[1] ^ phase_end[252][1]) || (phase_count[2] ^ phase_end[252][2]) || (phase_count[3] ^ phase_end[252][3]) || (phase_count[4] ^ phase_end[252][4]) || (phase_count[5] ^ phase_end[252][5]) || (phase_count[6] ^ phase_end[252][6]) || phase[252][7];
	assign select_end[253] = (phase_count[0] ^ phase_end[253][0]) || (phase_count[1] ^ phase_end[253][1]) || (phase_count[2] ^ phase_end[253][2]) || (phase_count[3] ^ phase_end[253][3]) || (phase_count[4] ^ phase_end[253][4]) || (phase_count[5] ^ phase_end[253][5]) || (phase_count[6] ^ phase_end[253][6]) || phase[253][7];
	assign select_end[254] = (phase_count[0] ^ phase_end[254][0]) || (phase_count[1] ^ phase_end[254][1]) || (phase_count[2] ^ phase_end[254][2]) || (phase_count[3] ^ phase_end[254][3]) || (phase_count[4] ^ phase_end[254][4]) || (phase_count[5] ^ phase_end[254][5]) || (phase_count[6] ^ phase_end[254][6]) || phase[254][7];
	assign select_end[255] = (phase_count[0] ^ phase_end[255][0]) || (phase_count[1] ^ phase_end[255][1]) || (phase_count[2] ^ phase_end[255][2]) || (phase_count[3] ^ phase_end[255][3]) || (phase_count[4] ^ phase_end[255][4]) || (phase_count[5] ^ phase_end[255][5]) || (phase_count[6] ^ phase_end[255][6]) || phase[255][7];
		
	//values is dependent on both the phase_clock and whether the select or select_end bits are 0;
	//assign values[0] = (values[0] & select[0] & select_end[0]) || ((phase_clock ^ (!((phase[0][5] & (phase[0][4] || phase[0][3])) || phase[0][6]))) & (!select[0]));
	//logic is as follows: values = itselft unless select or select_end are high. If select is high, value = 1. If select_end is high, value = 0;
	
	assign values[0] = (values[0] & select[0] & select_end[0]) || ((phase_clock ^ (!((phase[0][5] & (phase[0][4] || phase[0][3])) || phase[0][6]))) & (!select[0]));
	assign values[1] = (values[1] & select[1] & select_end[1]) || ((phase_clock ^ (!((phase[1][5] & (phase[1][4] || phase[1][3])) || phase[1][6]))) & (!select[1]));
	assign values[2] = (values[2] & select[2] & select_end[2]) || ((phase_clock ^ (!((phase[2][5] & (phase[2][4] || phase[2][3])) || phase[2][6]))) & (!select[2]));
	assign values[3] = (values[3] & select[3] & select_end[3]) || ((phase_clock ^ (!((phase[3][5] & (phase[3][4] || phase[3][3])) || phase[3][6]))) & (!select[3]));
	assign values[4] = (values[4] & select[4] & select_end[4]) || ((phase_clock ^ (!((phase[4][5] & (phase[4][4] || phase[4][3])) || phase[4][6]))) & (!select[4]));
	assign values[5] = (values[5] & select[5] & select_end[5]) || ((phase_clock ^ (!((phase[5][5] & (phase[5][4] || phase[5][3])) || phase[5][6]))) & (!select[5]));
	assign values[6] = (values[6] & select[6] & select_end[6]) || ((phase_clock ^ (!((phase[6][5] & (phase[6][4] || phase[6][3])) || phase[6][6]))) & (!select[6]));
	assign values[7] = (values[7] & select[7] & select_end[7]) || ((phase_clock ^ (!((phase[7][5] & (phase[7][4] || phase[7][3])) || phase[7][6]))) & (!select[7]));
	assign values[8] = (values[8] & select[8] & select_end[8]) || ((phase_clock ^ (!((phase[8][5] & (phase[8][4] || phase[8][3])) || phase[8][6]))) & (!select[8]));
	assign values[9] = (values[9] & select[9] & select_end[9]) || ((phase_clock ^ (!((phase[9][5] & (phase[9][4] || phase[9][3])) || phase[9][6]))) & (!select[9]));
	assign values[10] = (values[10] & select[10] & select_end[10]) || ((phase_clock ^ (!((phase[10][5] & (phase[10][4] || phase[10][3])) || phase[10][6]))) & (!select[10]));
	assign values[11] = (values[11] & select[11] & select_end[11]) || ((phase_clock ^ (!((phase[11][5] & (phase[11][4] || phase[11][3])) || phase[11][6]))) & (!select[11]));
	assign values[12] = (values[12] & select[12] & select_end[12]) || ((phase_clock ^ (!((phase[12][5] & (phase[12][4] || phase[12][3])) || phase[12][6]))) & (!select[12]));
	assign values[13] = (values[13] & select[13] & select_end[13]) || ((phase_clock ^ (!((phase[13][5] & (phase[13][4] || phase[13][3])) || phase[13][6]))) & (!select[13]));
	assign values[14] = (values[14] & select[14] & select_end[14]) || ((phase_clock ^ (!((phase[14][5] & (phase[14][4] || phase[14][3])) || phase[14][6]))) & (!select[14]));
	assign values[15] = (values[15] & select[15] & select_end[15]) || ((phase_clock ^ (!((phase[15][5] & (phase[15][4] || phase[15][3])) || phase[15][6]))) & (!select[15]));
	assign values[16] = (values[16] & select[16] & select_end[16]) || ((phase_clock ^ (!((phase[16][5] & (phase[16][4] || phase[16][3])) || phase[16][6]))) & (!select[16]));
	assign values[17] = (values[17] & select[17] & select_end[17]) || ((phase_clock ^ (!((phase[17][5] & (phase[17][4] || phase[17][3])) || phase[17][6]))) & (!select[17]));
	assign values[18] = (values[18] & select[18] & select_end[18]) || ((phase_clock ^ (!((phase[18][5] & (phase[18][4] || phase[18][3])) || phase[18][6]))) & (!select[18]));
	assign values[19] = (values[19] & select[19] & select_end[19]) || ((phase_clock ^ (!((phase[19][5] & (phase[19][4] || phase[19][3])) || phase[19][6]))) & (!select[19]));
	assign values[20] = (values[20] & select[20] & select_end[20]) || ((phase_clock ^ (!((phase[20][5] & (phase[20][4] || phase[20][3])) || phase[20][6]))) & (!select[20]));
	assign values[21] = (values[21] & select[21] & select_end[21]) || ((phase_clock ^ (!((phase[21][5] & (phase[21][4] || phase[21][3])) || phase[21][6]))) & (!select[21]));
	assign values[22] = (values[22] & select[22] & select_end[22]) || ((phase_clock ^ (!((phase[22][5] & (phase[22][4] || phase[22][3])) || phase[22][6]))) & (!select[22]));
	assign values[23] = (values[23] & select[23] & select_end[23]) || ((phase_clock ^ (!((phase[23][5] & (phase[23][4] || phase[23][3])) || phase[23][6]))) & (!select[23]));
	assign values[24] = (values[24] & select[24] & select_end[24]) || ((phase_clock ^ (!((phase[24][5] & (phase[24][4] || phase[24][3])) || phase[24][6]))) & (!select[24]));
	assign values[25] = (values[25] & select[25] & select_end[25]) || ((phase_clock ^ (!((phase[25][5] & (phase[25][4] || phase[25][3])) || phase[25][6]))) & (!select[25]));
	assign values[26] = (values[26] & select[26] & select_end[26]) || ((phase_clock ^ (!((phase[26][5] & (phase[26][4] || phase[26][3])) || phase[26][6]))) & (!select[26]));
	assign values[27] = (values[27] & select[27] & select_end[27]) || ((phase_clock ^ (!((phase[27][5] & (phase[27][4] || phase[27][3])) || phase[27][6]))) & (!select[27]));
	assign values[28] = (values[28] & select[28] & select_end[28]) || ((phase_clock ^ (!((phase[28][5] & (phase[28][4] || phase[28][3])) || phase[28][6]))) & (!select[28]));
	assign values[29] = (values[29] & select[29] & select_end[29]) || ((phase_clock ^ (!((phase[29][5] & (phase[29][4] || phase[29][3])) || phase[29][6]))) & (!select[29]));
	assign values[30] = (values[30] & select[30] & select_end[30]) || ((phase_clock ^ (!((phase[30][5] & (phase[30][4] || phase[30][3])) || phase[30][6]))) & (!select[30]));
	assign values[31] = (values[31] & select[31] & select_end[31]) || ((phase_clock ^ (!((phase[31][5] & (phase[31][4] || phase[31][3])) || phase[31][6]))) & (!select[31]));
	assign values[32] = (values[32] & select[32] & select_end[32]) || ((phase_clock ^ (!((phase[32][5] & (phase[32][4] || phase[32][3])) || phase[32][6]))) & (!select[32]));
	assign values[33] = (values[33] & select[33] & select_end[33]) || ((phase_clock ^ (!((phase[33][5] & (phase[33][4] || phase[33][3])) || phase[33][6]))) & (!select[33]));
	assign values[34] = (values[34] & select[34] & select_end[34]) || ((phase_clock ^ (!((phase[34][5] & (phase[34][4] || phase[34][3])) || phase[34][6]))) & (!select[34]));
	assign values[35] = (values[35] & select[35] & select_end[35]) || ((phase_clock ^ (!((phase[35][5] & (phase[35][4] || phase[35][3])) || phase[35][6]))) & (!select[35]));
	assign values[36] = (values[36] & select[36] & select_end[36]) || ((phase_clock ^ (!((phase[36][5] & (phase[36][4] || phase[36][3])) || phase[36][6]))) & (!select[36]));
	assign values[37] = (values[37] & select[37] & select_end[37]) || ((phase_clock ^ (!((phase[37][5] & (phase[37][4] || phase[37][3])) || phase[37][6]))) & (!select[37]));
	assign values[38] = (values[38] & select[38] & select_end[38]) || ((phase_clock ^ (!((phase[38][5] & (phase[38][4] || phase[38][3])) || phase[38][6]))) & (!select[38]));
	assign values[39] = (values[39] & select[39] & select_end[39]) || ((phase_clock ^ (!((phase[39][5] & (phase[39][4] || phase[39][3])) || phase[39][6]))) & (!select[39]));
	assign values[40] = (values[40] & select[40] & select_end[40]) || ((phase_clock ^ (!((phase[40][5] & (phase[40][4] || phase[40][3])) || phase[40][6]))) & (!select[40]));
	assign values[41] = (values[41] & select[41] & select_end[41]) || ((phase_clock ^ (!((phase[41][5] & (phase[41][4] || phase[41][3])) || phase[41][6]))) & (!select[41]));
	assign values[42] = (values[42] & select[42] & select_end[42]) || ((phase_clock ^ (!((phase[42][5] & (phase[42][4] || phase[42][3])) || phase[42][6]))) & (!select[42]));
	assign values[43] = (values[43] & select[43] & select_end[43]) || ((phase_clock ^ (!((phase[43][5] & (phase[43][4] || phase[43][3])) || phase[43][6]))) & (!select[43]));
	assign values[44] = (values[44] & select[44] & select_end[44]) || ((phase_clock ^ (!((phase[44][5] & (phase[44][4] || phase[44][3])) || phase[44][6]))) & (!select[44]));
	assign values[45] = (values[45] & select[45] & select_end[45]) || ((phase_clock ^ (!((phase[45][5] & (phase[45][4] || phase[45][3])) || phase[45][6]))) & (!select[45]));
	assign values[46] = (values[46] & select[46] & select_end[46]) || ((phase_clock ^ (!((phase[46][5] & (phase[46][4] || phase[46][3])) || phase[46][6]))) & (!select[46]));
	assign values[47] = (values[47] & select[47] & select_end[47]) || ((phase_clock ^ (!((phase[47][5] & (phase[47][4] || phase[47][3])) || phase[47][6]))) & (!select[47]));
	assign values[48] = (values[48] & select[48] & select_end[48]) || ((phase_clock ^ (!((phase[48][5] & (phase[48][4] || phase[48][3])) || phase[48][6]))) & (!select[48]));
	assign values[49] = (values[49] & select[49] & select_end[49]) || ((phase_clock ^ (!((phase[49][5] & (phase[49][4] || phase[49][3])) || phase[49][6]))) & (!select[49]));
	assign values[50] = (values[50] & select[50] & select_end[50]) || ((phase_clock ^ (!((phase[50][5] & (phase[50][4] || phase[50][3])) || phase[50][6]))) & (!select[50]));
	assign values[51] = (values[51] & select[51] & select_end[51]) || ((phase_clock ^ (!((phase[51][5] & (phase[51][4] || phase[51][3])) || phase[51][6]))) & (!select[51]));
	assign values[52] = (values[52] & select[52] & select_end[52]) || ((phase_clock ^ (!((phase[52][5] & (phase[52][4] || phase[52][3])) || phase[52][6]))) & (!select[52]));
	assign values[53] = (values[53] & select[53] & select_end[53]) || ((phase_clock ^ (!((phase[53][5] & (phase[53][4] || phase[53][3])) || phase[53][6]))) & (!select[53]));
	assign values[54] = (values[54] & select[54] & select_end[54]) || ((phase_clock ^ (!((phase[54][5] & (phase[54][4] || phase[54][3])) || phase[54][6]))) & (!select[54]));
	assign values[55] = (values[55] & select[55] & select_end[55]) || ((phase_clock ^ (!((phase[55][5] & (phase[55][4] || phase[55][3])) || phase[55][6]))) & (!select[55]));
	assign values[56] = (values[56] & select[56] & select_end[56]) || ((phase_clock ^ (!((phase[56][5] & (phase[56][4] || phase[56][3])) || phase[56][6]))) & (!select[56]));
	assign values[57] = (values[57] & select[57] & select_end[57]) || ((phase_clock ^ (!((phase[57][5] & (phase[57][4] || phase[57][3])) || phase[57][6]))) & (!select[57]));
	assign values[58] = (values[58] & select[58] & select_end[58]) || ((phase_clock ^ (!((phase[58][5] & (phase[58][4] || phase[58][3])) || phase[58][6]))) & (!select[58]));
	assign values[59] = (values[59] & select[59] & select_end[59]) || ((phase_clock ^ (!((phase[59][5] & (phase[59][4] || phase[59][3])) || phase[59][6]))) & (!select[59]));
	assign values[60] = (values[60] & select[60] & select_end[60]) || ((phase_clock ^ (!((phase[60][5] & (phase[60][4] || phase[60][3])) || phase[60][6]))) & (!select[60]));
	assign values[61] = (values[61] & select[61] & select_end[61]) || ((phase_clock ^ (!((phase[61][5] & (phase[61][4] || phase[61][3])) || phase[61][6]))) & (!select[61]));
	assign values[62] = (values[62] & select[62] & select_end[62]) || ((phase_clock ^ (!((phase[62][5] & (phase[62][4] || phase[62][3])) || phase[62][6]))) & (!select[62]));
	assign values[63] = (values[63] & select[63] & select_end[63]) || ((phase_clock ^ (!((phase[63][5] & (phase[63][4] || phase[63][3])) || phase[63][6]))) & (!select[63]));
	assign values[64] = (values[64] & select[64] & select_end[64]) || ((phase_clock ^ (!((phase[64][5] & (phase[64][4] || phase[64][3])) || phase[64][6]))) & (!select[64]));
	assign values[65] = (values[65] & select[65] & select_end[65]) || ((phase_clock ^ (!((phase[65][5] & (phase[65][4] || phase[65][3])) || phase[65][6]))) & (!select[65]));
	assign values[66] = (values[66] & select[66] & select_end[66]) || ((phase_clock ^ (!((phase[66][5] & (phase[66][4] || phase[66][3])) || phase[66][6]))) & (!select[66]));
	assign values[67] = (values[67] & select[67] & select_end[67]) || ((phase_clock ^ (!((phase[67][5] & (phase[67][4] || phase[67][3])) || phase[67][6]))) & (!select[67]));
	assign values[68] = (values[68] & select[68] & select_end[68]) || ((phase_clock ^ (!((phase[68][5] & (phase[68][4] || phase[68][3])) || phase[68][6]))) & (!select[68]));
	assign values[69] = (values[69] & select[69] & select_end[69]) || ((phase_clock ^ (!((phase[69][5] & (phase[69][4] || phase[69][3])) || phase[69][6]))) & (!select[69]));
	assign values[70] = (values[70] & select[70] & select_end[70]) || ((phase_clock ^ (!((phase[70][5] & (phase[70][4] || phase[70][3])) || phase[70][6]))) & (!select[70]));
	assign values[71] = (values[71] & select[71] & select_end[71]) || ((phase_clock ^ (!((phase[71][5] & (phase[71][4] || phase[71][3])) || phase[71][6]))) & (!select[71]));
	assign values[72] = (values[72] & select[72] & select_end[72]) || ((phase_clock ^ (!((phase[72][5] & (phase[72][4] || phase[72][3])) || phase[72][6]))) & (!select[72]));
	assign values[73] = (values[73] & select[73] & select_end[73]) || ((phase_clock ^ (!((phase[73][5] & (phase[73][4] || phase[73][3])) || phase[73][6]))) & (!select[73]));
	assign values[74] = (values[74] & select[74] & select_end[74]) || ((phase_clock ^ (!((phase[74][5] & (phase[74][4] || phase[74][3])) || phase[74][6]))) & (!select[74]));
	assign values[75] = (values[75] & select[75] & select_end[75]) || ((phase_clock ^ (!((phase[75][5] & (phase[75][4] || phase[75][3])) || phase[75][6]))) & (!select[75]));
	assign values[76] = (values[76] & select[76] & select_end[76]) || ((phase_clock ^ (!((phase[76][5] & (phase[76][4] || phase[76][3])) || phase[76][6]))) & (!select[76]));
	assign values[77] = (values[77] & select[77] & select_end[77]) || ((phase_clock ^ (!((phase[77][5] & (phase[77][4] || phase[77][3])) || phase[77][6]))) & (!select[77]));
	assign values[78] = (values[78] & select[78] & select_end[78]) || ((phase_clock ^ (!((phase[78][5] & (phase[78][4] || phase[78][3])) || phase[78][6]))) & (!select[78]));
	assign values[79] = (values[79] & select[79] & select_end[79]) || ((phase_clock ^ (!((phase[79][5] & (phase[79][4] || phase[79][3])) || phase[79][6]))) & (!select[79]));
	assign values[80] = (values[80] & select[80] & select_end[80]) || ((phase_clock ^ (!((phase[80][5] & (phase[80][4] || phase[80][3])) || phase[80][6]))) & (!select[80]));
	assign values[81] = (values[81] & select[81] & select_end[81]) || ((phase_clock ^ (!((phase[81][5] & (phase[81][4] || phase[81][3])) || phase[81][6]))) & (!select[81]));
	assign values[82] = (values[82] & select[82] & select_end[82]) || ((phase_clock ^ (!((phase[82][5] & (phase[82][4] || phase[82][3])) || phase[82][6]))) & (!select[82]));
	assign values[83] = (values[83] & select[83] & select_end[83]) || ((phase_clock ^ (!((phase[83][5] & (phase[83][4] || phase[83][3])) || phase[83][6]))) & (!select[83]));
	assign values[84] = (values[84] & select[84] & select_end[84]) || ((phase_clock ^ (!((phase[84][5] & (phase[84][4] || phase[84][3])) || phase[84][6]))) & (!select[84]));
	assign values[85] = (values[85] & select[85] & select_end[85]) || ((phase_clock ^ (!((phase[85][5] & (phase[85][4] || phase[85][3])) || phase[85][6]))) & (!select[85]));
	assign values[86] = (values[86] & select[86] & select_end[86]) || ((phase_clock ^ (!((phase[86][5] & (phase[86][4] || phase[86][3])) || phase[86][6]))) & (!select[86]));
	assign values[87] = (values[87] & select[87] & select_end[87]) || ((phase_clock ^ (!((phase[87][5] & (phase[87][4] || phase[87][3])) || phase[87][6]))) & (!select[87]));
	assign values[88] = (values[88] & select[88] & select_end[88]) || ((phase_clock ^ (!((phase[88][5] & (phase[88][4] || phase[88][3])) || phase[88][6]))) & (!select[88]));
	assign values[89] = (values[89] & select[89] & select_end[89]) || ((phase_clock ^ (!((phase[89][5] & (phase[89][4] || phase[89][3])) || phase[89][6]))) & (!select[89]));
	assign values[90] = (values[90] & select[90] & select_end[90]) || ((phase_clock ^ (!((phase[90][5] & (phase[90][4] || phase[90][3])) || phase[90][6]))) & (!select[90]));
	assign values[91] = (values[91] & select[91] & select_end[91]) || ((phase_clock ^ (!((phase[91][5] & (phase[91][4] || phase[91][3])) || phase[91][6]))) & (!select[91]));
	assign values[92] = (values[92] & select[92] & select_end[92]) || ((phase_clock ^ (!((phase[92][5] & (phase[92][4] || phase[92][3])) || phase[92][6]))) & (!select[92]));
	assign values[93] = (values[93] & select[93] & select_end[93]) || ((phase_clock ^ (!((phase[93][5] & (phase[93][4] || phase[93][3])) || phase[93][6]))) & (!select[93]));
	assign values[94] = (values[94] & select[94] & select_end[94]) || ((phase_clock ^ (!((phase[94][5] & (phase[94][4] || phase[94][3])) || phase[94][6]))) & (!select[94]));
	assign values[95] = (values[95] & select[95] & select_end[95]) || ((phase_clock ^ (!((phase[95][5] & (phase[95][4] || phase[95][3])) || phase[95][6]))) & (!select[95]));
	assign values[96] = (values[96] & select[96] & select_end[96]) || ((phase_clock ^ (!((phase[96][5] & (phase[96][4] || phase[96][3])) || phase[96][6]))) & (!select[96]));
	assign values[97] = (values[97] & select[97] & select_end[97]) || ((phase_clock ^ (!((phase[97][5] & (phase[97][4] || phase[97][3])) || phase[97][6]))) & (!select[97]));
	assign values[98] = (values[98] & select[98] & select_end[98]) || ((phase_clock ^ (!((phase[98][5] & (phase[98][4] || phase[98][3])) || phase[98][6]))) & (!select[98]));
	assign values[99] = (values[99] & select[99] & select_end[99]) || ((phase_clock ^ (!((phase[99][5] & (phase[99][4] || phase[99][3])) || phase[99][6]))) & (!select[99]));
	assign values[100] = (values[100] & select[100] & select_end[100]) || ((phase_clock ^ (!((phase[100][5] & (phase[100][4] || phase[100][3])) || phase[100][6]))) & (!select[100]));
	assign values[101] = (values[101] & select[101] & select_end[101]) || ((phase_clock ^ (!((phase[101][5] & (phase[101][4] || phase[101][3])) || phase[101][6]))) & (!select[101]));
	assign values[102] = (values[102] & select[102] & select_end[102]) || ((phase_clock ^ (!((phase[102][5] & (phase[102][4] || phase[102][3])) || phase[102][6]))) & (!select[102]));
	assign values[103] = (values[103] & select[103] & select_end[103]) || ((phase_clock ^ (!((phase[103][5] & (phase[103][4] || phase[103][3])) || phase[103][6]))) & (!select[103]));
	assign values[104] = (values[104] & select[104] & select_end[104]) || ((phase_clock ^ (!((phase[104][5] & (phase[104][4] || phase[104][3])) || phase[104][6]))) & (!select[104]));
	assign values[105] = (values[105] & select[105] & select_end[105]) || ((phase_clock ^ (!((phase[105][5] & (phase[105][4] || phase[105][3])) || phase[105][6]))) & (!select[105]));
	assign values[106] = (values[106] & select[106] & select_end[106]) || ((phase_clock ^ (!((phase[106][5] & (phase[106][4] || phase[106][3])) || phase[106][6]))) & (!select[106]));
	assign values[107] = (values[107] & select[107] & select_end[107]) || ((phase_clock ^ (!((phase[107][5] & (phase[107][4] || phase[107][3])) || phase[107][6]))) & (!select[107]));
	assign values[108] = (values[108] & select[108] & select_end[108]) || ((phase_clock ^ (!((phase[108][5] & (phase[108][4] || phase[108][3])) || phase[108][6]))) & (!select[108]));
	assign values[109] = (values[109] & select[109] & select_end[109]) || ((phase_clock ^ (!((phase[109][5] & (phase[109][4] || phase[109][3])) || phase[109][6]))) & (!select[109]));
	assign values[110] = (values[110] & select[110] & select_end[110]) || ((phase_clock ^ (!((phase[110][5] & (phase[110][4] || phase[110][3])) || phase[110][6]))) & (!select[110]));
	assign values[111] = (values[111] & select[111] & select_end[111]) || ((phase_clock ^ (!((phase[111][5] & (phase[111][4] || phase[111][3])) || phase[111][6]))) & (!select[111]));
	assign values[112] = (values[112] & select[112] & select_end[112]) || ((phase_clock ^ (!((phase[112][5] & (phase[112][4] || phase[112][3])) || phase[112][6]))) & (!select[112]));
	assign values[113] = (values[113] & select[113] & select_end[113]) || ((phase_clock ^ (!((phase[113][5] & (phase[113][4] || phase[113][3])) || phase[113][6]))) & (!select[113]));
	assign values[114] = (values[114] & select[114] & select_end[114]) || ((phase_clock ^ (!((phase[114][5] & (phase[114][4] || phase[114][3])) || phase[114][6]))) & (!select[114]));
	assign values[115] = (values[115] & select[115] & select_end[115]) || ((phase_clock ^ (!((phase[115][5] & (phase[115][4] || phase[115][3])) || phase[115][6]))) & (!select[115]));
	assign values[116] = (values[116] & select[116] & select_end[116]) || ((phase_clock ^ (!((phase[116][5] & (phase[116][4] || phase[116][3])) || phase[116][6]))) & (!select[116]));
	assign values[117] = (values[117] & select[117] & select_end[117]) || ((phase_clock ^ (!((phase[117][5] & (phase[117][4] || phase[117][3])) || phase[117][6]))) & (!select[117]));
	assign values[118] = (values[118] & select[118] & select_end[118]) || ((phase_clock ^ (!((phase[118][5] & (phase[118][4] || phase[118][3])) || phase[118][6]))) & (!select[118]));
	assign values[119] = (values[119] & select[119] & select_end[119]) || ((phase_clock ^ (!((phase[119][5] & (phase[119][4] || phase[119][3])) || phase[119][6]))) & (!select[119]));
	assign values[120] = (values[120] & select[120] & select_end[120]) || ((phase_clock ^ (!((phase[120][5] & (phase[120][4] || phase[120][3])) || phase[120][6]))) & (!select[120]));
	assign values[121] = (values[121] & select[121] & select_end[121]) || ((phase_clock ^ (!((phase[121][5] & (phase[121][4] || phase[121][3])) || phase[121][6]))) & (!select[121]));
	assign values[122] = (values[122] & select[122] & select_end[122]) || ((phase_clock ^ (!((phase[122][5] & (phase[122][4] || phase[122][3])) || phase[122][6]))) & (!select[122]));
	assign values[123] = (values[123] & select[123] & select_end[123]) || ((phase_clock ^ (!((phase[123][5] & (phase[123][4] || phase[123][3])) || phase[123][6]))) & (!select[123]));
	assign values[124] = (values[124] & select[124] & select_end[124]) || ((phase_clock ^ (!((phase[124][5] & (phase[124][4] || phase[124][3])) || phase[124][6]))) & (!select[124]));
	assign values[125] = (values[125] & select[125] & select_end[125]) || ((phase_clock ^ (!((phase[125][5] & (phase[125][4] || phase[125][3])) || phase[125][6]))) & (!select[125]));
	assign values[126] = (values[126] & select[126] & select_end[126]) || ((phase_clock ^ (!((phase[126][5] & (phase[126][4] || phase[126][3])) || phase[126][6]))) & (!select[126]));
	assign values[127] = (values[127] & select[127] & select_end[127]) || ((phase_clock ^ (!((phase[127][5] & (phase[127][4] || phase[127][3])) || phase[127][6]))) & (!select[127]));
	assign values[128] = (values[128] & select[128] & select_end[128]) || ((phase_clock ^ (!((phase[128][5] & (phase[128][4] || phase[128][3])) || phase[128][6]))) & (!select[128]));
	assign values[129] = (values[129] & select[129] & select_end[129]) || ((phase_clock ^ (!((phase[129][5] & (phase[129][4] || phase[129][3])) || phase[129][6]))) & (!select[129]));
	assign values[130] = (values[130] & select[130] & select_end[130]) || ((phase_clock ^ (!((phase[130][5] & (phase[130][4] || phase[130][3])) || phase[130][6]))) & (!select[130]));
	assign values[131] = (values[131] & select[131] & select_end[131]) || ((phase_clock ^ (!((phase[131][5] & (phase[131][4] || phase[131][3])) || phase[131][6]))) & (!select[131]));
	assign values[132] = (values[132] & select[132] & select_end[132]) || ((phase_clock ^ (!((phase[132][5] & (phase[132][4] || phase[132][3])) || phase[132][6]))) & (!select[132]));
	assign values[133] = (values[133] & select[133] & select_end[133]) || ((phase_clock ^ (!((phase[133][5] & (phase[133][4] || phase[133][3])) || phase[133][6]))) & (!select[133]));
	assign values[134] = (values[134] & select[134] & select_end[134]) || ((phase_clock ^ (!((phase[134][5] & (phase[134][4] || phase[134][3])) || phase[134][6]))) & (!select[134]));
	assign values[135] = (values[135] & select[135] & select_end[135]) || ((phase_clock ^ (!((phase[135][5] & (phase[135][4] || phase[135][3])) || phase[135][6]))) & (!select[135]));
	assign values[136] = (values[136] & select[136] & select_end[136]) || ((phase_clock ^ (!((phase[136][5] & (phase[136][4] || phase[136][3])) || phase[136][6]))) & (!select[136]));
	assign values[137] = (values[137] & select[137] & select_end[137]) || ((phase_clock ^ (!((phase[137][5] & (phase[137][4] || phase[137][3])) || phase[137][6]))) & (!select[137]));
	assign values[138] = (values[138] & select[138] & select_end[138]) || ((phase_clock ^ (!((phase[138][5] & (phase[138][4] || phase[138][3])) || phase[138][6]))) & (!select[138]));
	assign values[139] = (values[139] & select[139] & select_end[139]) || ((phase_clock ^ (!((phase[139][5] & (phase[139][4] || phase[139][3])) || phase[139][6]))) & (!select[139]));
	assign values[140] = (values[140] & select[140] & select_end[140]) || ((phase_clock ^ (!((phase[140][5] & (phase[140][4] || phase[140][3])) || phase[140][6]))) & (!select[140]));
	assign values[141] = (values[141] & select[141] & select_end[141]) || ((phase_clock ^ (!((phase[141][5] & (phase[141][4] || phase[141][3])) || phase[141][6]))) & (!select[141]));
	assign values[142] = (values[142] & select[142] & select_end[142]) || ((phase_clock ^ (!((phase[142][5] & (phase[142][4] || phase[142][3])) || phase[142][6]))) & (!select[142]));
	assign values[143] = (values[143] & select[143] & select_end[143]) || ((phase_clock ^ (!((phase[143][5] & (phase[143][4] || phase[143][3])) || phase[143][6]))) & (!select[143]));
	assign values[144] = (values[144] & select[144] & select_end[144]) || ((phase_clock ^ (!((phase[144][5] & (phase[144][4] || phase[144][3])) || phase[144][6]))) & (!select[144]));
	assign values[145] = (values[145] & select[145] & select_end[145]) || ((phase_clock ^ (!((phase[145][5] & (phase[145][4] || phase[145][3])) || phase[145][6]))) & (!select[145]));
	assign values[146] = (values[146] & select[146] & select_end[146]) || ((phase_clock ^ (!((phase[146][5] & (phase[146][4] || phase[146][3])) || phase[146][6]))) & (!select[146]));
	assign values[147] = (values[147] & select[147] & select_end[147]) || ((phase_clock ^ (!((phase[147][5] & (phase[147][4] || phase[147][3])) || phase[147][6]))) & (!select[147]));
	assign values[148] = (values[148] & select[148] & select_end[148]) || ((phase_clock ^ (!((phase[148][5] & (phase[148][4] || phase[148][3])) || phase[148][6]))) & (!select[148]));
	assign values[149] = (values[149] & select[149] & select_end[149]) || ((phase_clock ^ (!((phase[149][5] & (phase[149][4] || phase[149][3])) || phase[149][6]))) & (!select[149]));
	assign values[150] = (values[150] & select[150] & select_end[150]) || ((phase_clock ^ (!((phase[150][5] & (phase[150][4] || phase[150][3])) || phase[150][6]))) & (!select[150]));
	assign values[151] = (values[151] & select[151] & select_end[151]) || ((phase_clock ^ (!((phase[151][5] & (phase[151][4] || phase[151][3])) || phase[151][6]))) & (!select[151]));
	assign values[152] = (values[152] & select[152] & select_end[152]) || ((phase_clock ^ (!((phase[152][5] & (phase[152][4] || phase[152][3])) || phase[152][6]))) & (!select[152]));
	assign values[153] = (values[153] & select[153] & select_end[153]) || ((phase_clock ^ (!((phase[153][5] & (phase[153][4] || phase[153][3])) || phase[153][6]))) & (!select[153]));
	assign values[154] = (values[154] & select[154] & select_end[154]) || ((phase_clock ^ (!((phase[154][5] & (phase[154][4] || phase[154][3])) || phase[154][6]))) & (!select[154]));
	assign values[155] = (values[155] & select[155] & select_end[155]) || ((phase_clock ^ (!((phase[155][5] & (phase[155][4] || phase[155][3])) || phase[155][6]))) & (!select[155]));
	assign values[156] = (values[156] & select[156] & select_end[156]) || ((phase_clock ^ (!((phase[156][5] & (phase[156][4] || phase[156][3])) || phase[156][6]))) & (!select[156]));
	assign values[157] = (values[157] & select[157] & select_end[157]) || ((phase_clock ^ (!((phase[157][5] & (phase[157][4] || phase[157][3])) || phase[157][6]))) & (!select[157]));
	assign values[158] = (values[158] & select[158] & select_end[158]) || ((phase_clock ^ (!((phase[158][5] & (phase[158][4] || phase[158][3])) || phase[158][6]))) & (!select[158]));
	assign values[159] = (values[159] & select[159] & select_end[159]) || ((phase_clock ^ (!((phase[159][5] & (phase[159][4] || phase[159][3])) || phase[159][6]))) & (!select[159]));
	assign values[160] = (values[160] & select[160] & select_end[160]) || ((phase_clock ^ (!((phase[160][5] & (phase[160][4] || phase[160][3])) || phase[160][6]))) & (!select[160]));
	assign values[161] = (values[161] & select[161] & select_end[161]) || ((phase_clock ^ (!((phase[161][5] & (phase[161][4] || phase[161][3])) || phase[161][6]))) & (!select[161]));
	assign values[162] = (values[162] & select[162] & select_end[162]) || ((phase_clock ^ (!((phase[162][5] & (phase[162][4] || phase[162][3])) || phase[162][6]))) & (!select[162]));
	assign values[163] = (values[163] & select[163] & select_end[163]) || ((phase_clock ^ (!((phase[163][5] & (phase[163][4] || phase[163][3])) || phase[163][6]))) & (!select[163]));
	assign values[164] = (values[164] & select[164] & select_end[164]) || ((phase_clock ^ (!((phase[164][5] & (phase[164][4] || phase[164][3])) || phase[164][6]))) & (!select[164]));
	assign values[165] = (values[165] & select[165] & select_end[165]) || ((phase_clock ^ (!((phase[165][5] & (phase[165][4] || phase[165][3])) || phase[165][6]))) & (!select[165]));
	assign values[166] = (values[166] & select[166] & select_end[166]) || ((phase_clock ^ (!((phase[166][5] & (phase[166][4] || phase[166][3])) || phase[166][6]))) & (!select[166]));
	assign values[167] = (values[167] & select[167] & select_end[167]) || ((phase_clock ^ (!((phase[167][5] & (phase[167][4] || phase[167][3])) || phase[167][6]))) & (!select[167]));
	assign values[168] = (values[168] & select[168] & select_end[168]) || ((phase_clock ^ (!((phase[168][5] & (phase[168][4] || phase[168][3])) || phase[168][6]))) & (!select[168]));
	assign values[169] = (values[169] & select[169] & select_end[169]) || ((phase_clock ^ (!((phase[169][5] & (phase[169][4] || phase[169][3])) || phase[169][6]))) & (!select[169]));
	assign values[170] = (values[170] & select[170] & select_end[170]) || ((phase_clock ^ (!((phase[170][5] & (phase[170][4] || phase[170][3])) || phase[170][6]))) & (!select[170]));
	assign values[171] = (values[171] & select[171] & select_end[171]) || ((phase_clock ^ (!((phase[171][5] & (phase[171][4] || phase[171][3])) || phase[171][6]))) & (!select[171]));
	assign values[172] = (values[172] & select[172] & select_end[172]) || ((phase_clock ^ (!((phase[172][5] & (phase[172][4] || phase[172][3])) || phase[172][6]))) & (!select[172]));
	assign values[173] = (values[173] & select[173] & select_end[173]) || ((phase_clock ^ (!((phase[173][5] & (phase[173][4] || phase[173][3])) || phase[173][6]))) & (!select[173]));
	assign values[174] = (values[174] & select[174] & select_end[174]) || ((phase_clock ^ (!((phase[174][5] & (phase[174][4] || phase[174][3])) || phase[174][6]))) & (!select[174]));
	assign values[175] = (values[175] & select[175] & select_end[175]) || ((phase_clock ^ (!((phase[175][5] & (phase[175][4] || phase[175][3])) || phase[175][6]))) & (!select[175]));
	assign values[176] = (values[176] & select[176] & select_end[176]) || ((phase_clock ^ (!((phase[176][5] & (phase[176][4] || phase[176][3])) || phase[176][6]))) & (!select[176]));
	assign values[177] = (values[177] & select[177] & select_end[177]) || ((phase_clock ^ (!((phase[177][5] & (phase[177][4] || phase[177][3])) || phase[177][6]))) & (!select[177]));
	assign values[178] = (values[178] & select[178] & select_end[178]) || ((phase_clock ^ (!((phase[178][5] & (phase[178][4] || phase[178][3])) || phase[178][6]))) & (!select[178]));
	assign values[179] = (values[179] & select[179] & select_end[179]) || ((phase_clock ^ (!((phase[179][5] & (phase[179][4] || phase[179][3])) || phase[179][6]))) & (!select[179]));
	assign values[180] = (values[180] & select[180] & select_end[180]) || ((phase_clock ^ (!((phase[180][5] & (phase[180][4] || phase[180][3])) || phase[180][6]))) & (!select[180]));
	assign values[181] = (values[181] & select[181] & select_end[181]) || ((phase_clock ^ (!((phase[181][5] & (phase[181][4] || phase[181][3])) || phase[181][6]))) & (!select[181]));
	assign values[182] = (values[182] & select[182] & select_end[182]) || ((phase_clock ^ (!((phase[182][5] & (phase[182][4] || phase[182][3])) || phase[182][6]))) & (!select[182]));
	assign values[183] = (values[183] & select[183] & select_end[183]) || ((phase_clock ^ (!((phase[183][5] & (phase[183][4] || phase[183][3])) || phase[183][6]))) & (!select[183]));
	assign values[184] = (values[184] & select[184] & select_end[184]) || ((phase_clock ^ (!((phase[184][5] & (phase[184][4] || phase[184][3])) || phase[184][6]))) & (!select[184]));
	assign values[185] = (values[185] & select[185] & select_end[185]) || ((phase_clock ^ (!((phase[185][5] & (phase[185][4] || phase[185][3])) || phase[185][6]))) & (!select[185]));
	assign values[186] = (values[186] & select[186] & select_end[186]) || ((phase_clock ^ (!((phase[186][5] & (phase[186][4] || phase[186][3])) || phase[186][6]))) & (!select[186]));
	assign values[187] = (values[187] & select[187] & select_end[187]) || ((phase_clock ^ (!((phase[187][5] & (phase[187][4] || phase[187][3])) || phase[187][6]))) & (!select[187]));
	assign values[188] = (values[188] & select[188] & select_end[188]) || ((phase_clock ^ (!((phase[188][5] & (phase[188][4] || phase[188][3])) || phase[188][6]))) & (!select[188]));
	assign values[189] = (values[189] & select[189] & select_end[189]) || ((phase_clock ^ (!((phase[189][5] & (phase[189][4] || phase[189][3])) || phase[189][6]))) & (!select[189]));
	assign values[190] = (values[190] & select[190] & select_end[190]) || ((phase_clock ^ (!((phase[190][5] & (phase[190][4] || phase[190][3])) || phase[190][6]))) & (!select[190]));
	assign values[191] = (values[191] & select[191] & select_end[191]) || ((phase_clock ^ (!((phase[191][5] & (phase[191][4] || phase[191][3])) || phase[191][6]))) & (!select[191]));
	assign values[192] = (values[192] & select[192] & select_end[192]) || ((phase_clock ^ (!((phase[192][5] & (phase[192][4] || phase[192][3])) || phase[192][6]))) & (!select[192]));
	assign values[193] = (values[193] & select[193] & select_end[193]) || ((phase_clock ^ (!((phase[193][5] & (phase[193][4] || phase[193][3])) || phase[193][6]))) & (!select[193]));
	assign values[194] = (values[194] & select[194] & select_end[194]) || ((phase_clock ^ (!((phase[194][5] & (phase[194][4] || phase[194][3])) || phase[194][6]))) & (!select[194]));
	assign values[195] = (values[195] & select[195] & select_end[195]) || ((phase_clock ^ (!((phase[195][5] & (phase[195][4] || phase[195][3])) || phase[195][6]))) & (!select[195]));
	assign values[196] = (values[196] & select[196] & select_end[196]) || ((phase_clock ^ (!((phase[196][5] & (phase[196][4] || phase[196][3])) || phase[196][6]))) & (!select[196]));
	assign values[197] = (values[197] & select[197] & select_end[197]) || ((phase_clock ^ (!((phase[197][5] & (phase[197][4] || phase[197][3])) || phase[197][6]))) & (!select[197]));
	assign values[198] = (values[198] & select[198] & select_end[198]) || ((phase_clock ^ (!((phase[198][5] & (phase[198][4] || phase[198][3])) || phase[198][6]))) & (!select[198]));
	assign values[199] = (values[199] & select[199] & select_end[199]) || ((phase_clock ^ (!((phase[199][5] & (phase[199][4] || phase[199][3])) || phase[199][6]))) & (!select[199]));
	assign values[200] = (values[200] & select[200] & select_end[200]) || ((phase_clock ^ (!((phase[200][5] & (phase[200][4] || phase[200][3])) || phase[200][6]))) & (!select[200]));
	assign values[201] = (values[201] & select[201] & select_end[201]) || ((phase_clock ^ (!((phase[201][5] & (phase[201][4] || phase[201][3])) || phase[201][6]))) & (!select[201]));
	assign values[202] = (values[202] & select[202] & select_end[202]) || ((phase_clock ^ (!((phase[202][5] & (phase[202][4] || phase[202][3])) || phase[202][6]))) & (!select[202]));
	assign values[203] = (values[203] & select[203] & select_end[203]) || ((phase_clock ^ (!((phase[203][5] & (phase[203][4] || phase[203][3])) || phase[203][6]))) & (!select[203]));
	assign values[204] = (values[204] & select[204] & select_end[204]) || ((phase_clock ^ (!((phase[204][5] & (phase[204][4] || phase[204][3])) || phase[204][6]))) & (!select[204]));
	assign values[205] = (values[205] & select[205] & select_end[205]) || ((phase_clock ^ (!((phase[205][5] & (phase[205][4] || phase[205][3])) || phase[205][6]))) & (!select[205]));
	assign values[206] = (values[206] & select[206] & select_end[206]) || ((phase_clock ^ (!((phase[206][5] & (phase[206][4] || phase[206][3])) || phase[206][6]))) & (!select[206]));
	assign values[207] = (values[207] & select[207] & select_end[207]) || ((phase_clock ^ (!((phase[207][5] & (phase[207][4] || phase[207][3])) || phase[207][6]))) & (!select[207]));
	assign values[208] = (values[208] & select[208] & select_end[208]) || ((phase_clock ^ (!((phase[208][5] & (phase[208][4] || phase[208][3])) || phase[208][6]))) & (!select[208]));
	assign values[209] = (values[209] & select[209] & select_end[209]) || ((phase_clock ^ (!((phase[209][5] & (phase[209][4] || phase[209][3])) || phase[209][6]))) & (!select[209]));
	assign values[210] = (values[210] & select[210] & select_end[210]) || ((phase_clock ^ (!((phase[210][5] & (phase[210][4] || phase[210][3])) || phase[210][6]))) & (!select[210]));
	assign values[211] = (values[211] & select[211] & select_end[211]) || ((phase_clock ^ (!((phase[211][5] & (phase[211][4] || phase[211][3])) || phase[211][6]))) & (!select[211]));
	assign values[212] = (values[212] & select[212] & select_end[212]) || ((phase_clock ^ (!((phase[212][5] & (phase[212][4] || phase[212][3])) || phase[212][6]))) & (!select[212]));
	assign values[213] = (values[213] & select[213] & select_end[213]) || ((phase_clock ^ (!((phase[213][5] & (phase[213][4] || phase[213][3])) || phase[213][6]))) & (!select[213]));
	assign values[214] = (values[214] & select[214] & select_end[214]) || ((phase_clock ^ (!((phase[214][5] & (phase[214][4] || phase[214][3])) || phase[214][6]))) & (!select[214]));
	assign values[215] = (values[215] & select[215] & select_end[215]) || ((phase_clock ^ (!((phase[215][5] & (phase[215][4] || phase[215][3])) || phase[215][6]))) & (!select[215]));
	assign values[216] = (values[216] & select[216] & select_end[216]) || ((phase_clock ^ (!((phase[216][5] & (phase[216][4] || phase[216][3])) || phase[216][6]))) & (!select[216]));
	assign values[217] = (values[217] & select[217] & select_end[217]) || ((phase_clock ^ (!((phase[217][5] & (phase[217][4] || phase[217][3])) || phase[217][6]))) & (!select[217]));
	assign values[218] = (values[218] & select[218] & select_end[218]) || ((phase_clock ^ (!((phase[218][5] & (phase[218][4] || phase[218][3])) || phase[218][6]))) & (!select[218]));
	assign values[219] = (values[219] & select[219] & select_end[219]) || ((phase_clock ^ (!((phase[219][5] & (phase[219][4] || phase[219][3])) || phase[219][6]))) & (!select[219]));
	assign values[220] = (values[220] & select[220] & select_end[220]) || ((phase_clock ^ (!((phase[220][5] & (phase[220][4] || phase[220][3])) || phase[220][6]))) & (!select[220]));
	assign values[221] = (values[221] & select[221] & select_end[221]) || ((phase_clock ^ (!((phase[221][5] & (phase[221][4] || phase[221][3])) || phase[221][6]))) & (!select[221]));
	assign values[222] = (values[222] & select[222] & select_end[222]) || ((phase_clock ^ (!((phase[222][5] & (phase[222][4] || phase[222][3])) || phase[222][6]))) & (!select[222]));
	assign values[223] = (values[223] & select[223] & select_end[223]) || ((phase_clock ^ (!((phase[223][5] & (phase[223][4] || phase[223][3])) || phase[223][6]))) & (!select[223]));
	assign values[224] = (values[224] & select[224] & select_end[224]) || ((phase_clock ^ (!((phase[224][5] & (phase[224][4] || phase[224][3])) || phase[224][6]))) & (!select[224]));
	assign values[225] = (values[225] & select[225] & select_end[225]) || ((phase_clock ^ (!((phase[225][5] & (phase[225][4] || phase[225][3])) || phase[225][6]))) & (!select[225]));
	assign values[226] = (values[226] & select[226] & select_end[226]) || ((phase_clock ^ (!((phase[226][5] & (phase[226][4] || phase[226][3])) || phase[226][6]))) & (!select[226]));
	assign values[227] = (values[227] & select[227] & select_end[227]) || ((phase_clock ^ (!((phase[227][5] & (phase[227][4] || phase[227][3])) || phase[227][6]))) & (!select[227]));
	assign values[228] = (values[228] & select[228] & select_end[228]) || ((phase_clock ^ (!((phase[228][5] & (phase[228][4] || phase[228][3])) || phase[228][6]))) & (!select[228]));
	assign values[229] = (values[229] & select[229] & select_end[229]) || ((phase_clock ^ (!((phase[229][5] & (phase[229][4] || phase[229][3])) || phase[229][6]))) & (!select[229]));
	assign values[230] = (values[230] & select[230] & select_end[230]) || ((phase_clock ^ (!((phase[230][5] & (phase[230][4] || phase[230][3])) || phase[230][6]))) & (!select[230]));
	assign values[231] = (values[231] & select[231] & select_end[231]) || ((phase_clock ^ (!((phase[231][5] & (phase[231][4] || phase[231][3])) || phase[231][6]))) & (!select[231]));
	assign values[232] = (values[232] & select[232] & select_end[232]) || ((phase_clock ^ (!((phase[232][5] & (phase[232][4] || phase[232][3])) || phase[232][6]))) & (!select[232]));
	assign values[233] = (values[233] & select[233] & select_end[233]) || ((phase_clock ^ (!((phase[233][5] & (phase[233][4] || phase[233][3])) || phase[233][6]))) & (!select[233]));
	assign values[234] = (values[234] & select[234] & select_end[234]) || ((phase_clock ^ (!((phase[234][5] & (phase[234][4] || phase[234][3])) || phase[234][6]))) & (!select[234]));
	assign values[235] = (values[235] & select[235] & select_end[235]) || ((phase_clock ^ (!((phase[235][5] & (phase[235][4] || phase[235][3])) || phase[235][6]))) & (!select[235]));
	assign values[236] = (values[236] & select[236] & select_end[236]) || ((phase_clock ^ (!((phase[236][5] & (phase[236][4] || phase[236][3])) || phase[236][6]))) & (!select[236]));
	assign values[237] = (values[237] & select[237] & select_end[237]) || ((phase_clock ^ (!((phase[237][5] & (phase[237][4] || phase[237][3])) || phase[237][6]))) & (!select[237]));
	assign values[238] = (values[238] & select[238] & select_end[238]) || ((phase_clock ^ (!((phase[238][5] & (phase[238][4] || phase[238][3])) || phase[238][6]))) & (!select[238]));
	assign values[239] = (values[239] & select[239] & select_end[239]) || ((phase_clock ^ (!((phase[239][5] & (phase[239][4] || phase[239][3])) || phase[239][6]))) & (!select[239]));
	assign values[240] = (values[240] & select[240] & select_end[240]) || ((phase_clock ^ (!((phase[240][5] & (phase[240][4] || phase[240][3])) || phase[240][6]))) & (!select[240]));
	assign values[241] = (values[241] & select[241] & select_end[241]) || ((phase_clock ^ (!((phase[241][5] & (phase[241][4] || phase[241][3])) || phase[241][6]))) & (!select[241]));
	assign values[242] = (values[242] & select[242] & select_end[242]) || ((phase_clock ^ (!((phase[242][5] & (phase[242][4] || phase[242][3])) || phase[242][6]))) & (!select[242]));
	assign values[243] = (values[243] & select[243] & select_end[243]) || ((phase_clock ^ (!((phase[243][5] & (phase[243][4] || phase[243][3])) || phase[243][6]))) & (!select[243]));
	assign values[244] = (values[244] & select[244] & select_end[244]) || ((phase_clock ^ (!((phase[244][5] & (phase[244][4] || phase[244][3])) || phase[244][6]))) & (!select[244]));
	assign values[245] = (values[245] & select[245] & select_end[245]) || ((phase_clock ^ (!((phase[245][5] & (phase[245][4] || phase[245][3])) || phase[245][6]))) & (!select[245]));
	assign values[246] = (values[246] & select[246] & select_end[246]) || ((phase_clock ^ (!((phase[246][5] & (phase[246][4] || phase[246][3])) || phase[246][6]))) & (!select[246]));
	assign values[247] = (values[247] & select[247] & select_end[247]) || ((phase_clock ^ (!((phase[247][5] & (phase[247][4] || phase[247][3])) || phase[247][6]))) & (!select[247]));
	assign values[248] = (values[248] & select[248] & select_end[248]) || ((phase_clock ^ (!((phase[248][5] & (phase[248][4] || phase[248][3])) || phase[248][6]))) & (!select[248]));
	assign values[249] = (values[249] & select[249] & select_end[249]) || ((phase_clock ^ (!((phase[249][5] & (phase[249][4] || phase[249][3])) || phase[249][6]))) & (!select[249]));
	assign values[250] = (values[250] & select[250] & select_end[250]) || ((phase_clock ^ (!((phase[250][5] & (phase[250][4] || phase[250][3])) || phase[250][6]))) & (!select[250]));
	assign values[251] = (values[251] & select[251] & select_end[251]) || ((phase_clock ^ (!((phase[251][5] & (phase[251][4] || phase[251][3])) || phase[251][6]))) & (!select[251]));
	assign values[252] = (values[252] & select[252] & select_end[252]) || ((phase_clock ^ (!((phase[252][5] & (phase[252][4] || phase[252][3])) || phase[252][6]))) & (!select[252]));
	assign values[253] = (values[253] & select[253] & select_end[253]) || ((phase_clock ^ (!((phase[253][5] & (phase[253][4] || phase[253][3])) || phase[253][6]))) & (!select[253]));
	assign values[254] = (values[254] & select[254] & select_end[254]) || ((phase_clock ^ (!((phase[254][5] & (phase[254][4] || phase[254][3])) || phase[254][6]))) & (!select[254]));
	assign values[255] = (values[255] & select[255] & select_end[255]) || ((phase_clock ^ (!((phase[255][5] & (phase[255][4] || phase[255][3])) || phase[255][6]))) & (!select[255]));
			
	//output bits in order 32 bits at a time
	assign dataOut[0] = values[0 + counter[2:0]] & cnt[17];
	assign dataOut[1] = values[8 + counter[2:0]] & cnt[17];
	assign dataOut[2] = values[16 + counter[2:0]] & cnt[17];
	assign dataOut[3] = values[24 + counter[2:0]] & cnt[17];
	assign dataOut[4] = values[32 + counter[2:0]] & cnt[17];
	assign dataOut[5] = values[40 + counter[2:0]] & cnt[17];
	assign dataOut[6] = values[48 + counter[2:0]] & cnt[17];
	assign dataOut[7] = values[56 + counter[2:0]] & cnt[17];
	assign dataOut[8] = values[64 + counter[2:0]] & cnt[17];
	assign dataOut[9] = values[72 + counter[2:0]] & cnt[17];
	assign dataOut[10] = values[80 + counter[2:0]] & cnt[17];
	assign dataOut[11] = values[88 + counter[2:0]] & cnt[17];
	assign dataOut[12] = values[96 + counter[2:0]] & cnt[17];
	assign dataOut[13] = values[104 + counter[2:0]] & cnt[17];
	assign dataOut[14] = values[112 + counter[2:0]] & cnt[17];
	assign dataOut[15] = values[120 + counter[2:0]] & cnt[17];
	assign dataOut[16] = values[128 + counter[2:0]] & cnt[17];
	assign dataOut[17] = values[136 + counter[2:0]] & cnt[17];
	assign dataOut[18] = values[144 + counter[2:0]] & cnt[17];
	assign dataOut[19] = values[152 + counter[2:0]] & cnt[17];
	assign dataOut[20] = values[160 + counter[2:0]] & cnt[17];
	assign dataOut[21] = values[168 + counter[2:0]] & cnt[17];
	assign dataOut[22] = values[176 + counter[2:0]] & cnt[17];
	assign dataOut[23] = values[184 + counter[2:0]] & cnt[17];
	assign dataOut[24] = values[192 + counter[2:0]] & cnt[17];
	assign dataOut[25] = values[200 + counter[2:0]] & cnt[17];
	assign dataOut[26] = values[208 + counter[2:0]] & cnt[17];
	assign dataOut[27] = values[216 + counter[2:0]] & cnt[17];
	assign dataOut[28] = values[224 + counter[2:0]] & cnt[17];
	assign dataOut[29] = values[232 + counter[2:0]] & cnt[17];
	assign dataOut[30] = values[240 + counter[2:0]] & cnt[17];
	assign dataOut[31] = values[248 + counter[2:0]] & cnt[17];
	
	//testing pin
	assign clkOut = cnt[0];
	//the latch gate is 1/32 the speed of the normal clock
	assign latch = !(cnt[0] || cnt[1] || cnt[2] || cnt[3]);
	//each latch clock covers half the PCB
	assign latch2 = !(cnt[0] || cnt[1] || cnt[2] || cnt[3]);
	//take two input uart clocks at the same speed with slight offset and xor them to make a faster clock to read uart input
	assign uart_clock = uart_clock1 ^ uart_clock2;
	//testing pin
	assign clkCompare2 = uart_clock;

endmodule
