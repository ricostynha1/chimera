// This program was cloned from: https://github.com/scalabletoeplitz/HDL-Bits
// License: The Unlicense

module top_module(
    output zero
);// Module body starts after semicolon

    assign zero = 2'b00;
    
endmodule
