// This program was cloned from: https://github.com/Nilesh002/Multiplication-and-Accumulation-Unit-MAC-
// License: MIT License

module add48(a,b,s);
input [47:0]a,b;
output [47:0]s;

assign s=a+b;

endmodule
