// This program was cloned from: https://github.com/WangXuan95/FPGA-Gzip-compressor
// License: GNU General Public License v3.0


module static_huffman_table (
    input  wire        clk,
    input  wire [ 8:0] i_symbol,
    output wire [ 8:0] o_huffman_bits,
    output wire [ 3:0] o_huffman_len
);

reg  [ 8:0] bits;
reg  [ 3:0] len;

assign o_huffman_bits = bits;
assign o_huffman_len  = len;

always @ (posedge clk)
    case (i_symbol)
        9'h000 : begin  bits <= 9'h00c;  len <= 4'd8;  end
        9'h001 : begin  bits <= 9'h08c;  len <= 4'd8;  end
        9'h002 : begin  bits <= 9'h04c;  len <= 4'd8;  end
        9'h003 : begin  bits <= 9'h0cc;  len <= 4'd8;  end
        9'h004 : begin  bits <= 9'h02c;  len <= 4'd8;  end
        9'h005 : begin  bits <= 9'h0ac;  len <= 4'd8;  end
        9'h006 : begin  bits <= 9'h06c;  len <= 4'd8;  end
        9'h007 : begin  bits <= 9'h0ec;  len <= 4'd8;  end
        9'h008 : begin  bits <= 9'h01c;  len <= 4'd8;  end
        9'h009 : begin  bits <= 9'h09c;  len <= 4'd8;  end
        9'h00a : begin  bits <= 9'h05c;  len <= 4'd8;  end
        9'h00b : begin  bits <= 9'h0dc;  len <= 4'd8;  end
        9'h00c : begin  bits <= 9'h03c;  len <= 4'd8;  end
        9'h00d : begin  bits <= 9'h0bc;  len <= 4'd8;  end
        9'h00e : begin  bits <= 9'h07c;  len <= 4'd8;  end
        9'h00f : begin  bits <= 9'h0fc;  len <= 4'd8;  end
        9'h010 : begin  bits <= 9'h002;  len <= 4'd8;  end
        9'h011 : begin  bits <= 9'h082;  len <= 4'd8;  end
        9'h012 : begin  bits <= 9'h042;  len <= 4'd8;  end
        9'h013 : begin  bits <= 9'h0c2;  len <= 4'd8;  end
        9'h014 : begin  bits <= 9'h022;  len <= 4'd8;  end
        9'h015 : begin  bits <= 9'h0a2;  len <= 4'd8;  end
        9'h016 : begin  bits <= 9'h062;  len <= 4'd8;  end
        9'h017 : begin  bits <= 9'h0e2;  len <= 4'd8;  end
        9'h018 : begin  bits <= 9'h012;  len <= 4'd8;  end
        9'h019 : begin  bits <= 9'h092;  len <= 4'd8;  end
        9'h01a : begin  bits <= 9'h052;  len <= 4'd8;  end
        9'h01b : begin  bits <= 9'h0d2;  len <= 4'd8;  end
        9'h01c : begin  bits <= 9'h032;  len <= 4'd8;  end
        9'h01d : begin  bits <= 9'h0b2;  len <= 4'd8;  end
        9'h01e : begin  bits <= 9'h072;  len <= 4'd8;  end
        9'h01f : begin  bits <= 9'h0f2;  len <= 4'd8;  end
        9'h020 : begin  bits <= 9'h00a;  len <= 4'd8;  end
        9'h021 : begin  bits <= 9'h08a;  len <= 4'd8;  end
        9'h022 : begin  bits <= 9'h04a;  len <= 4'd8;  end
        9'h023 : begin  bits <= 9'h0ca;  len <= 4'd8;  end
        9'h024 : begin  bits <= 9'h02a;  len <= 4'd8;  end
        9'h025 : begin  bits <= 9'h0aa;  len <= 4'd8;  end
        9'h026 : begin  bits <= 9'h06a;  len <= 4'd8;  end
        9'h027 : begin  bits <= 9'h0ea;  len <= 4'd8;  end
        9'h028 : begin  bits <= 9'h01a;  len <= 4'd8;  end
        9'h029 : begin  bits <= 9'h09a;  len <= 4'd8;  end
        9'h02a : begin  bits <= 9'h05a;  len <= 4'd8;  end
        9'h02b : begin  bits <= 9'h0da;  len <= 4'd8;  end
        9'h02c : begin  bits <= 9'h03a;  len <= 4'd8;  end
        9'h02d : begin  bits <= 9'h0ba;  len <= 4'd8;  end
        9'h02e : begin  bits <= 9'h07a;  len <= 4'd8;  end
        9'h02f : begin  bits <= 9'h0fa;  len <= 4'd8;  end
        9'h030 : begin  bits <= 9'h006;  len <= 4'd8;  end
        9'h031 : begin  bits <= 9'h086;  len <= 4'd8;  end
        9'h032 : begin  bits <= 9'h046;  len <= 4'd8;  end
        9'h033 : begin  bits <= 9'h0c6;  len <= 4'd8;  end
        9'h034 : begin  bits <= 9'h026;  len <= 4'd8;  end
        9'h035 : begin  bits <= 9'h0a6;  len <= 4'd8;  end
        9'h036 : begin  bits <= 9'h066;  len <= 4'd8;  end
        9'h037 : begin  bits <= 9'h0e6;  len <= 4'd8;  end
        9'h038 : begin  bits <= 9'h016;  len <= 4'd8;  end
        9'h039 : begin  bits <= 9'h096;  len <= 4'd8;  end
        9'h03a : begin  bits <= 9'h056;  len <= 4'd8;  end
        9'h03b : begin  bits <= 9'h0d6;  len <= 4'd8;  end
        9'h03c : begin  bits <= 9'h036;  len <= 4'd8;  end
        9'h03d : begin  bits <= 9'h0b6;  len <= 4'd8;  end
        9'h03e : begin  bits <= 9'h076;  len <= 4'd8;  end
        9'h03f : begin  bits <= 9'h0f6;  len <= 4'd8;  end
        9'h040 : begin  bits <= 9'h00e;  len <= 4'd8;  end
        9'h041 : begin  bits <= 9'h08e;  len <= 4'd8;  end
        9'h042 : begin  bits <= 9'h04e;  len <= 4'd8;  end
        9'h043 : begin  bits <= 9'h0ce;  len <= 4'd8;  end
        9'h044 : begin  bits <= 9'h02e;  len <= 4'd8;  end
        9'h045 : begin  bits <= 9'h0ae;  len <= 4'd8;  end
        9'h046 : begin  bits <= 9'h06e;  len <= 4'd8;  end
        9'h047 : begin  bits <= 9'h0ee;  len <= 4'd8;  end
        9'h048 : begin  bits <= 9'h01e;  len <= 4'd8;  end
        9'h049 : begin  bits <= 9'h09e;  len <= 4'd8;  end
        9'h04a : begin  bits <= 9'h05e;  len <= 4'd8;  end
        9'h04b : begin  bits <= 9'h0de;  len <= 4'd8;  end
        9'h04c : begin  bits <= 9'h03e;  len <= 4'd8;  end
        9'h04d : begin  bits <= 9'h0be;  len <= 4'd8;  end
        9'h04e : begin  bits <= 9'h07e;  len <= 4'd8;  end
        9'h04f : begin  bits <= 9'h0fe;  len <= 4'd8;  end
        9'h050 : begin  bits <= 9'h001;  len <= 4'd8;  end
        9'h051 : begin  bits <= 9'h081;  len <= 4'd8;  end
        9'h052 : begin  bits <= 9'h041;  len <= 4'd8;  end
        9'h053 : begin  bits <= 9'h0c1;  len <= 4'd8;  end
        9'h054 : begin  bits <= 9'h021;  len <= 4'd8;  end
        9'h055 : begin  bits <= 9'h0a1;  len <= 4'd8;  end
        9'h056 : begin  bits <= 9'h061;  len <= 4'd8;  end
        9'h057 : begin  bits <= 9'h0e1;  len <= 4'd8;  end
        9'h058 : begin  bits <= 9'h011;  len <= 4'd8;  end
        9'h059 : begin  bits <= 9'h091;  len <= 4'd8;  end
        9'h05a : begin  bits <= 9'h051;  len <= 4'd8;  end
        9'h05b : begin  bits <= 9'h0d1;  len <= 4'd8;  end
        9'h05c : begin  bits <= 9'h031;  len <= 4'd8;  end
        9'h05d : begin  bits <= 9'h0b1;  len <= 4'd8;  end
        9'h05e : begin  bits <= 9'h071;  len <= 4'd8;  end
        9'h05f : begin  bits <= 9'h0f1;  len <= 4'd8;  end
        9'h060 : begin  bits <= 9'h009;  len <= 4'd8;  end
        9'h061 : begin  bits <= 9'h089;  len <= 4'd8;  end
        9'h062 : begin  bits <= 9'h049;  len <= 4'd8;  end
        9'h063 : begin  bits <= 9'h0c9;  len <= 4'd8;  end
        9'h064 : begin  bits <= 9'h029;  len <= 4'd8;  end
        9'h065 : begin  bits <= 9'h0a9;  len <= 4'd8;  end
        9'h066 : begin  bits <= 9'h069;  len <= 4'd8;  end
        9'h067 : begin  bits <= 9'h0e9;  len <= 4'd8;  end
        9'h068 : begin  bits <= 9'h019;  len <= 4'd8;  end
        9'h069 : begin  bits <= 9'h099;  len <= 4'd8;  end
        9'h06a : begin  bits <= 9'h059;  len <= 4'd8;  end
        9'h06b : begin  bits <= 9'h0d9;  len <= 4'd8;  end
        9'h06c : begin  bits <= 9'h039;  len <= 4'd8;  end
        9'h06d : begin  bits <= 9'h0b9;  len <= 4'd8;  end
        9'h06e : begin  bits <= 9'h079;  len <= 4'd8;  end
        9'h06f : begin  bits <= 9'h0f9;  len <= 4'd8;  end
        9'h070 : begin  bits <= 9'h005;  len <= 4'd8;  end
        9'h071 : begin  bits <= 9'h085;  len <= 4'd8;  end
        9'h072 : begin  bits <= 9'h045;  len <= 4'd8;  end
        9'h073 : begin  bits <= 9'h0c5;  len <= 4'd8;  end
        9'h074 : begin  bits <= 9'h025;  len <= 4'd8;  end
        9'h075 : begin  bits <= 9'h0a5;  len <= 4'd8;  end
        9'h076 : begin  bits <= 9'h065;  len <= 4'd8;  end
        9'h077 : begin  bits <= 9'h0e5;  len <= 4'd8;  end
        9'h078 : begin  bits <= 9'h015;  len <= 4'd8;  end
        9'h079 : begin  bits <= 9'h095;  len <= 4'd8;  end
        9'h07a : begin  bits <= 9'h055;  len <= 4'd8;  end
        9'h07b : begin  bits <= 9'h0d5;  len <= 4'd8;  end
        9'h07c : begin  bits <= 9'h035;  len <= 4'd8;  end
        9'h07d : begin  bits <= 9'h0b5;  len <= 4'd8;  end
        9'h07e : begin  bits <= 9'h075;  len <= 4'd8;  end
        9'h07f : begin  bits <= 9'h0f5;  len <= 4'd8;  end
        9'h080 : begin  bits <= 9'h00d;  len <= 4'd8;  end
        9'h081 : begin  bits <= 9'h08d;  len <= 4'd8;  end
        9'h082 : begin  bits <= 9'h04d;  len <= 4'd8;  end
        9'h083 : begin  bits <= 9'h0cd;  len <= 4'd8;  end
        9'h084 : begin  bits <= 9'h02d;  len <= 4'd8;  end
        9'h085 : begin  bits <= 9'h0ad;  len <= 4'd8;  end
        9'h086 : begin  bits <= 9'h06d;  len <= 4'd8;  end
        9'h087 : begin  bits <= 9'h0ed;  len <= 4'd8;  end
        9'h088 : begin  bits <= 9'h01d;  len <= 4'd8;  end
        9'h089 : begin  bits <= 9'h09d;  len <= 4'd8;  end
        9'h08a : begin  bits <= 9'h05d;  len <= 4'd8;  end
        9'h08b : begin  bits <= 9'h0dd;  len <= 4'd8;  end
        9'h08c : begin  bits <= 9'h03d;  len <= 4'd8;  end
        9'h08d : begin  bits <= 9'h0bd;  len <= 4'd8;  end
        9'h08e : begin  bits <= 9'h07d;  len <= 4'd8;  end
        9'h08f : begin  bits <= 9'h0fd;  len <= 4'd8;  end
        9'h090 : begin  bits <= 9'h013;  len <= 4'd9;  end
        9'h091 : begin  bits <= 9'h113;  len <= 4'd9;  end
        9'h092 : begin  bits <= 9'h093;  len <= 4'd9;  end
        9'h093 : begin  bits <= 9'h193;  len <= 4'd9;  end
        9'h094 : begin  bits <= 9'h053;  len <= 4'd9;  end
        9'h095 : begin  bits <= 9'h153;  len <= 4'd9;  end
        9'h096 : begin  bits <= 9'h0d3;  len <= 4'd9;  end
        9'h097 : begin  bits <= 9'h1d3;  len <= 4'd9;  end
        9'h098 : begin  bits <= 9'h033;  len <= 4'd9;  end
        9'h099 : begin  bits <= 9'h133;  len <= 4'd9;  end
        9'h09a : begin  bits <= 9'h0b3;  len <= 4'd9;  end
        9'h09b : begin  bits <= 9'h1b3;  len <= 4'd9;  end
        9'h09c : begin  bits <= 9'h073;  len <= 4'd9;  end
        9'h09d : begin  bits <= 9'h173;  len <= 4'd9;  end
        9'h09e : begin  bits <= 9'h0f3;  len <= 4'd9;  end
        9'h09f : begin  bits <= 9'h1f3;  len <= 4'd9;  end
        9'h0a0 : begin  bits <= 9'h00b;  len <= 4'd9;  end
        9'h0a1 : begin  bits <= 9'h10b;  len <= 4'd9;  end
        9'h0a2 : begin  bits <= 9'h08b;  len <= 4'd9;  end
        9'h0a3 : begin  bits <= 9'h18b;  len <= 4'd9;  end
        9'h0a4 : begin  bits <= 9'h04b;  len <= 4'd9;  end
        9'h0a5 : begin  bits <= 9'h14b;  len <= 4'd9;  end
        9'h0a6 : begin  bits <= 9'h0cb;  len <= 4'd9;  end
        9'h0a7 : begin  bits <= 9'h1cb;  len <= 4'd9;  end
        9'h0a8 : begin  bits <= 9'h02b;  len <= 4'd9;  end
        9'h0a9 : begin  bits <= 9'h12b;  len <= 4'd9;  end
        9'h0aa : begin  bits <= 9'h0ab;  len <= 4'd9;  end
        9'h0ab : begin  bits <= 9'h1ab;  len <= 4'd9;  end
        9'h0ac : begin  bits <= 9'h06b;  len <= 4'd9;  end
        9'h0ad : begin  bits <= 9'h16b;  len <= 4'd9;  end
        9'h0ae : begin  bits <= 9'h0eb;  len <= 4'd9;  end
        9'h0af : begin  bits <= 9'h1eb;  len <= 4'd9;  end
        9'h0b0 : begin  bits <= 9'h01b;  len <= 4'd9;  end
        9'h0b1 : begin  bits <= 9'h11b;  len <= 4'd9;  end
        9'h0b2 : begin  bits <= 9'h09b;  len <= 4'd9;  end
        9'h0b3 : begin  bits <= 9'h19b;  len <= 4'd9;  end
        9'h0b4 : begin  bits <= 9'h05b;  len <= 4'd9;  end
        9'h0b5 : begin  bits <= 9'h15b;  len <= 4'd9;  end
        9'h0b6 : begin  bits <= 9'h0db;  len <= 4'd9;  end
        9'h0b7 : begin  bits <= 9'h1db;  len <= 4'd9;  end
        9'h0b8 : begin  bits <= 9'h03b;  len <= 4'd9;  end
        9'h0b9 : begin  bits <= 9'h13b;  len <= 4'd9;  end
        9'h0ba : begin  bits <= 9'h0bb;  len <= 4'd9;  end
        9'h0bb : begin  bits <= 9'h1bb;  len <= 4'd9;  end
        9'h0bc : begin  bits <= 9'h07b;  len <= 4'd9;  end
        9'h0bd : begin  bits <= 9'h17b;  len <= 4'd9;  end
        9'h0be : begin  bits <= 9'h0fb;  len <= 4'd9;  end
        9'h0bf : begin  bits <= 9'h1fb;  len <= 4'd9;  end
        9'h0c0 : begin  bits <= 9'h007;  len <= 4'd9;  end
        9'h0c1 : begin  bits <= 9'h107;  len <= 4'd9;  end
        9'h0c2 : begin  bits <= 9'h087;  len <= 4'd9;  end
        9'h0c3 : begin  bits <= 9'h187;  len <= 4'd9;  end
        9'h0c4 : begin  bits <= 9'h047;  len <= 4'd9;  end
        9'h0c5 : begin  bits <= 9'h147;  len <= 4'd9;  end
        9'h0c6 : begin  bits <= 9'h0c7;  len <= 4'd9;  end
        9'h0c7 : begin  bits <= 9'h1c7;  len <= 4'd9;  end
        9'h0c8 : begin  bits <= 9'h027;  len <= 4'd9;  end
        9'h0c9 : begin  bits <= 9'h127;  len <= 4'd9;  end
        9'h0ca : begin  bits <= 9'h0a7;  len <= 4'd9;  end
        9'h0cb : begin  bits <= 9'h1a7;  len <= 4'd9;  end
        9'h0cc : begin  bits <= 9'h067;  len <= 4'd9;  end
        9'h0cd : begin  bits <= 9'h167;  len <= 4'd9;  end
        9'h0ce : begin  bits <= 9'h0e7;  len <= 4'd9;  end
        9'h0cf : begin  bits <= 9'h1e7;  len <= 4'd9;  end
        9'h0d0 : begin  bits <= 9'h017;  len <= 4'd9;  end
        9'h0d1 : begin  bits <= 9'h117;  len <= 4'd9;  end
        9'h0d2 : begin  bits <= 9'h097;  len <= 4'd9;  end
        9'h0d3 : begin  bits <= 9'h197;  len <= 4'd9;  end
        9'h0d4 : begin  bits <= 9'h057;  len <= 4'd9;  end
        9'h0d5 : begin  bits <= 9'h157;  len <= 4'd9;  end
        9'h0d6 : begin  bits <= 9'h0d7;  len <= 4'd9;  end
        9'h0d7 : begin  bits <= 9'h1d7;  len <= 4'd9;  end
        9'h0d8 : begin  bits <= 9'h037;  len <= 4'd9;  end
        9'h0d9 : begin  bits <= 9'h137;  len <= 4'd9;  end
        9'h0da : begin  bits <= 9'h0b7;  len <= 4'd9;  end
        9'h0db : begin  bits <= 9'h1b7;  len <= 4'd9;  end
        9'h0dc : begin  bits <= 9'h077;  len <= 4'd9;  end
        9'h0dd : begin  bits <= 9'h177;  len <= 4'd9;  end
        9'h0de : begin  bits <= 9'h0f7;  len <= 4'd9;  end
        9'h0df : begin  bits <= 9'h1f7;  len <= 4'd9;  end
        9'h0e0 : begin  bits <= 9'h00f;  len <= 4'd9;  end
        9'h0e1 : begin  bits <= 9'h10f;  len <= 4'd9;  end
        9'h0e2 : begin  bits <= 9'h08f;  len <= 4'd9;  end
        9'h0e3 : begin  bits <= 9'h18f;  len <= 4'd9;  end
        9'h0e4 : begin  bits <= 9'h04f;  len <= 4'd9;  end
        9'h0e5 : begin  bits <= 9'h14f;  len <= 4'd9;  end
        9'h0e6 : begin  bits <= 9'h0cf;  len <= 4'd9;  end
        9'h0e7 : begin  bits <= 9'h1cf;  len <= 4'd9;  end
        9'h0e8 : begin  bits <= 9'h02f;  len <= 4'd9;  end
        9'h0e9 : begin  bits <= 9'h12f;  len <= 4'd9;  end
        9'h0ea : begin  bits <= 9'h0af;  len <= 4'd9;  end
        9'h0eb : begin  bits <= 9'h1af;  len <= 4'd9;  end
        9'h0ec : begin  bits <= 9'h06f;  len <= 4'd9;  end
        9'h0ed : begin  bits <= 9'h16f;  len <= 4'd9;  end
        9'h0ee : begin  bits <= 9'h0ef;  len <= 4'd9;  end
        9'h0ef : begin  bits <= 9'h1ef;  len <= 4'd9;  end
        9'h0f0 : begin  bits <= 9'h01f;  len <= 4'd9;  end
        9'h0f1 : begin  bits <= 9'h11f;  len <= 4'd9;  end
        9'h0f2 : begin  bits <= 9'h09f;  len <= 4'd9;  end
        9'h0f3 : begin  bits <= 9'h19f;  len <= 4'd9;  end
        9'h0f4 : begin  bits <= 9'h05f;  len <= 4'd9;  end
        9'h0f5 : begin  bits <= 9'h15f;  len <= 4'd9;  end
        9'h0f6 : begin  bits <= 9'h0df;  len <= 4'd9;  end
        9'h0f7 : begin  bits <= 9'h1df;  len <= 4'd9;  end
        9'h0f8 : begin  bits <= 9'h03f;  len <= 4'd9;  end
        9'h0f9 : begin  bits <= 9'h13f;  len <= 4'd9;  end
        9'h0fa : begin  bits <= 9'h0bf;  len <= 4'd9;  end
        9'h0fb : begin  bits <= 9'h1bf;  len <= 4'd9;  end
        9'h0fc : begin  bits <= 9'h07f;  len <= 4'd9;  end
        9'h0fd : begin  bits <= 9'h17f;  len <= 4'd9;  end
        9'h0fe : begin  bits <= 9'h0ff;  len <= 4'd9;  end
        9'h0ff : begin  bits <= 9'h1ff;  len <= 4'd9;  end
        9'h100 : begin  bits <= 9'h000;  len <= 4'd7;  end
        9'h101 : begin  bits <= 9'h040;  len <= 4'd7;  end
        9'h102 : begin  bits <= 9'h020;  len <= 4'd7;  end
        9'h103 : begin  bits <= 9'h060;  len <= 4'd7;  end
        9'h104 : begin  bits <= 9'h010;  len <= 4'd7;  end
        9'h105 : begin  bits <= 9'h050;  len <= 4'd7;  end
        9'h106 : begin  bits <= 9'h030;  len <= 4'd7;  end
        9'h107 : begin  bits <= 9'h070;  len <= 4'd7;  end
        9'h108 : begin  bits <= 9'h008;  len <= 4'd7;  end
        9'h109 : begin  bits <= 9'h048;  len <= 4'd7;  end
        9'h10a : begin  bits <= 9'h028;  len <= 4'd7;  end
        9'h10b : begin  bits <= 9'h068;  len <= 4'd7;  end
        9'h10c : begin  bits <= 9'h018;  len <= 4'd7;  end
        9'h10d : begin  bits <= 9'h058;  len <= 4'd7;  end
        9'h10e : begin  bits <= 9'h038;  len <= 4'd7;  end
        9'h10f : begin  bits <= 9'h078;  len <= 4'd7;  end
        9'h110 : begin  bits <= 9'h004;  len <= 4'd7;  end
        9'h111 : begin  bits <= 9'h044;  len <= 4'd7;  end
        9'h112 : begin  bits <= 9'h024;  len <= 4'd7;  end
        9'h113 : begin  bits <= 9'h064;  len <= 4'd7;  end
        9'h114 : begin  bits <= 9'h014;  len <= 4'd7;  end
        9'h115 : begin  bits <= 9'h054;  len <= 4'd7;  end
        9'h116 : begin  bits <= 9'h034;  len <= 4'd7;  end
        9'h117 : begin  bits <= 9'h074;  len <= 4'd7;  end
        9'h118 : begin  bits <= 9'h003;  len <= 4'd8;  end
        9'h119 : begin  bits <= 9'h083;  len <= 4'd8;  end
        9'h11a : begin  bits <= 9'h043;  len <= 4'd8;  end
        9'h11b : begin  bits <= 9'h0c3;  len <= 4'd8;  end
        9'h11c : begin  bits <= 9'h023;  len <= 4'd8;  end
        9'h11d : begin  bits <= 9'h0a3;  len <= 4'd8;  end
        default: begin  bits <= 9'h0;    len <= 4'd0;  end
    endcase

endmodule
