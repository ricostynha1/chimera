// This program was cloned from: https://github.com/apuder/TRS-IO
// License: GNU General Public License v3.0

`timescale 1ns / 1ps

module videodetector(
   input vgaclk, // 25.2MHz clock
   input hsync_in,
   input vsync_in,

   output reg present,
   output reg hertz50
);


// Detect if the video input is present by measuring the period of the
// horizontal sync.  If it toggles with approximately the correct period
// then declare video as present.
// Detect if the video input is 60Hz or 50Hz by counting the number of
// horizontal scan rows.  Compare to the value midway between the number
// for 60 and 50 and if less than declare as 60Hz and if greater declare
// as 50Hz.
 
reg [1:0] hsync_in_dly;
reg [1:0] vsync_in_dly;

always @ (posedge vgaclk)
begin
   hsync_in_dly <= { hsync_in_dly[0], hsync_in }; // no glitch suppression
   //hsync_in_dly <= { hsync_in_dly[0], (^hsync_in_dly) ? hsync_in_dly[0] : hsync_in }; // glitch suppression

   vsync_in_dly[0] <= vsync_in; // no glitch suppression
end


// The horizontal rate is 15.84kHz.  25.2MHz/15.84kHz = 1591
reg [10:0] hcnt; // mod 1591 horizontal counter -1590..0 when hsync present

// The vertical rate is either 60Hz or 50Hz.  The 60Hz has 22 character rows,
// the 50Hz has 26 character rows.  Each character row is 12 scan rows.
// Detect 60/50 Hz by counting the scan rows per frame using a threshold of
// 24*12 = 288.
reg [8:0] vcnt;

always @ (posedge vgaclk)
begin
   // When present the hsync will sample xcnt when it crosses through zero.
   // The hsync signal is generated by a one-shot so only one edge is reliable
   // which from observation is the rising edge.
   if(hsync_in_dly == 2'b01) // rising edge
   begin
      // If the hsync is in the neighborhood of zero crossing then indicate
      // that video is present.
      present <= (hcnt[10:5] == 6'b111111 || hcnt[10:5] == 6'b000000) ? 1'b1: 1'b0;
      hcnt <= -11'd1590;

      vsync_in_dly[1] <= vsync_in_dly[0];
      if(vsync_in_dly == 2'b10) // falling edge
      begin
         hertz50 <= ~vcnt[8];
         vcnt <= -9'd287;
      end
      else
         vcnt <= vcnt + 9'd1;
   end
   else
   begin
      hcnt <= hcnt + 11'd1;
      // If counter wraps then must be free-running (no sync) so indicate
      // that video is not present.
      if(hcnt == -11'd1591)
         present <= 1'b0;
   end
end

endmodule
